VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu
  CLASS BLOCK ;
  FOREIGN alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN AluA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 39.480 350.000 40.080 ;
    END
  END AluA[0]
  PIN AluA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 66.680 350.000 67.280 ;
    END
  END AluA[10]
  PIN AluA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 69.400 350.000 70.000 ;
    END
  END AluA[11]
  PIN AluA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 72.120 350.000 72.720 ;
    END
  END AluA[12]
  PIN AluA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 74.840 350.000 75.440 ;
    END
  END AluA[13]
  PIN AluA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 77.560 350.000 78.160 ;
    END
  END AluA[14]
  PIN AluA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 80.280 350.000 80.880 ;
    END
  END AluA[15]
  PIN AluA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 83.000 350.000 83.600 ;
    END
  END AluA[16]
  PIN AluA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 85.720 350.000 86.320 ;
    END
  END AluA[17]
  PIN AluA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 88.440 350.000 89.040 ;
    END
  END AluA[18]
  PIN AluA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 91.160 350.000 91.760 ;
    END
  END AluA[19]
  PIN AluA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 42.200 350.000 42.800 ;
    END
  END AluA[1]
  PIN AluA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 93.880 350.000 94.480 ;
    END
  END AluA[20]
  PIN AluA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 96.600 350.000 97.200 ;
    END
  END AluA[21]
  PIN AluA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 346.000 99.320 350.000 99.920 ;
    END
  END AluA[22]
  PIN AluA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 102.040 350.000 102.640 ;
    END
  END AluA[23]
  PIN AluA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 104.760 350.000 105.360 ;
    END
  END AluA[24]
  PIN AluA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 107.480 350.000 108.080 ;
    END
  END AluA[25]
  PIN AluA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 346.000 110.200 350.000 110.800 ;
    END
  END AluA[26]
  PIN AluA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 112.920 350.000 113.520 ;
    END
  END AluA[27]
  PIN AluA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 115.640 350.000 116.240 ;
    END
  END AluA[28]
  PIN AluA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 118.360 350.000 118.960 ;
    END
  END AluA[29]
  PIN AluA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 44.920 350.000 45.520 ;
    END
  END AluA[2]
  PIN AluA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 121.080 350.000 121.680 ;
    END
  END AluA[30]
  PIN AluA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 123.800 350.000 124.400 ;
    END
  END AluA[31]
  PIN AluA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 47.640 350.000 48.240 ;
    END
  END AluA[3]
  PIN AluA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 50.360 350.000 50.960 ;
    END
  END AluA[4]
  PIN AluA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 53.080 350.000 53.680 ;
    END
  END AluA[5]
  PIN AluA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 55.800 350.000 56.400 ;
    END
  END AluA[6]
  PIN AluA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 58.520 350.000 59.120 ;
    END
  END AluA[7]
  PIN AluA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 61.240 350.000 61.840 ;
    END
  END AluA[8]
  PIN AluA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 63.960 350.000 64.560 ;
    END
  END AluA[9]
  PIN AluB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 126.520 350.000 127.120 ;
    END
  END AluB[0]
  PIN AluB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 153.720 350.000 154.320 ;
    END
  END AluB[10]
  PIN AluB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 156.440 350.000 157.040 ;
    END
  END AluB[11]
  PIN AluB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 159.160 350.000 159.760 ;
    END
  END AluB[12]
  PIN AluB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 161.880 350.000 162.480 ;
    END
  END AluB[13]
  PIN AluB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 164.600 350.000 165.200 ;
    END
  END AluB[14]
  PIN AluB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 167.320 350.000 167.920 ;
    END
  END AluB[15]
  PIN AluB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 170.040 350.000 170.640 ;
    END
  END AluB[16]
  PIN AluB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 172.760 350.000 173.360 ;
    END
  END AluB[17]
  PIN AluB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 175.480 350.000 176.080 ;
    END
  END AluB[18]
  PIN AluB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 178.200 350.000 178.800 ;
    END
  END AluB[19]
  PIN AluB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 129.240 350.000 129.840 ;
    END
  END AluB[1]
  PIN AluB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 180.920 350.000 181.520 ;
    END
  END AluB[20]
  PIN AluB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 183.640 350.000 184.240 ;
    END
  END AluB[21]
  PIN AluB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 186.360 350.000 186.960 ;
    END
  END AluB[22]
  PIN AluB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 189.080 350.000 189.680 ;
    END
  END AluB[23]
  PIN AluB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 191.800 350.000 192.400 ;
    END
  END AluB[24]
  PIN AluB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 194.520 350.000 195.120 ;
    END
  END AluB[25]
  PIN AluB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 197.240 350.000 197.840 ;
    END
  END AluB[26]
  PIN AluB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 199.960 350.000 200.560 ;
    END
  END AluB[27]
  PIN AluB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 202.680 350.000 203.280 ;
    END
  END AluB[28]
  PIN AluB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 205.400 350.000 206.000 ;
    END
  END AluB[29]
  PIN AluB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 131.960 350.000 132.560 ;
    END
  END AluB[2]
  PIN AluB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 208.120 350.000 208.720 ;
    END
  END AluB[30]
  PIN AluB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 210.840 350.000 211.440 ;
    END
  END AluB[31]
  PIN AluB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 134.680 350.000 135.280 ;
    END
  END AluB[3]
  PIN AluB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 137.400 350.000 138.000 ;
    END
  END AluB[4]
  PIN AluB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 140.120 350.000 140.720 ;
    END
  END AluB[5]
  PIN AluB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 142.840 350.000 143.440 ;
    END
  END AluB[6]
  PIN AluB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 145.560 350.000 146.160 ;
    END
  END AluB[7]
  PIN AluB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 148.280 350.000 148.880 ;
    END
  END AluB[8]
  PIN AluB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 151.000 350.000 151.600 ;
    END
  END AluB[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END VPWR
  PIN alucontrol[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 213.560 350.000 214.160 ;
    END
  END alucontrol[0]
  PIN alucontrol[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 216.280 350.000 216.880 ;
    END
  END alucontrol[1]
  PIN alucontrol[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 219.000 350.000 219.600 ;
    END
  END alucontrol[2]
  PIN alucontrol[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 221.720 350.000 222.320 ;
    END
  END alucontrol[3]
  PIN alucontrol[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 224.440 350.000 225.040 ;
    END
  END alucontrol[4]
  PIN aludone
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 227.160 350.000 227.760 ;
    END
  END aludone
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 346.000 34.040 350.000 34.640 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 36.760 350.000 37.360 ;
    END
  END reset
  PIN result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 229.880 350.000 230.480 ;
    END
  END result[0]
  PIN result[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 257.080 350.000 257.680 ;
    END
  END result[10]
  PIN result[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 259.800 350.000 260.400 ;
    END
  END result[11]
  PIN result[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 262.520 350.000 263.120 ;
    END
  END result[12]
  PIN result[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 265.240 350.000 265.840 ;
    END
  END result[13]
  PIN result[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 267.960 350.000 268.560 ;
    END
  END result[14]
  PIN result[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 270.680 350.000 271.280 ;
    END
  END result[15]
  PIN result[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 273.400 350.000 274.000 ;
    END
  END result[16]
  PIN result[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 276.120 350.000 276.720 ;
    END
  END result[17]
  PIN result[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 278.840 350.000 279.440 ;
    END
  END result[18]
  PIN result[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 281.560 350.000 282.160 ;
    END
  END result[19]
  PIN result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 232.600 350.000 233.200 ;
    END
  END result[1]
  PIN result[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 284.280 350.000 284.880 ;
    END
  END result[20]
  PIN result[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 287.000 350.000 287.600 ;
    END
  END result[21]
  PIN result[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 289.720 350.000 290.320 ;
    END
  END result[22]
  PIN result[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 292.440 350.000 293.040 ;
    END
  END result[23]
  PIN result[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 295.160 350.000 295.760 ;
    END
  END result[24]
  PIN result[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 297.880 350.000 298.480 ;
    END
  END result[25]
  PIN result[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 300.600 350.000 301.200 ;
    END
  END result[26]
  PIN result[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 303.320 350.000 303.920 ;
    END
  END result[27]
  PIN result[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 306.040 350.000 306.640 ;
    END
  END result[28]
  PIN result[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 308.760 350.000 309.360 ;
    END
  END result[29]
  PIN result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 235.320 350.000 235.920 ;
    END
  END result[2]
  PIN result[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 311.480 350.000 312.080 ;
    END
  END result[30]
  PIN result[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 314.200 350.000 314.800 ;
    END
  END result[31]
  PIN result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 238.040 350.000 238.640 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 240.760 350.000 241.360 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 243.480 350.000 244.080 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 246.200 350.000 246.800 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 248.920 350.000 249.520 ;
    END
  END result[7]
  PIN result[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 346.000 251.640 350.000 252.240 ;
    END
  END result[8]
  PIN result[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 346.000 254.360 350.000 254.960 ;
    END
  END result[9]
  OBS
      LAYER nwell ;
        RECT 5.330 333.145 344.270 335.975 ;
        RECT 5.330 327.705 344.270 330.535 ;
        RECT 5.330 322.265 344.270 325.095 ;
        RECT 5.330 316.825 344.270 319.655 ;
        RECT 5.330 311.385 344.270 314.215 ;
        RECT 5.330 305.945 344.270 308.775 ;
        RECT 5.330 300.505 344.270 303.335 ;
        RECT 5.330 295.065 344.270 297.895 ;
        RECT 5.330 289.625 344.270 292.455 ;
        RECT 5.330 284.185 344.270 287.015 ;
        RECT 5.330 278.745 344.270 281.575 ;
        RECT 5.330 273.305 344.270 276.135 ;
        RECT 5.330 267.865 344.270 270.695 ;
        RECT 5.330 262.425 344.270 265.255 ;
        RECT 5.330 256.985 344.270 259.815 ;
        RECT 5.330 251.545 344.270 254.375 ;
        RECT 5.330 246.105 344.270 248.935 ;
        RECT 5.330 240.665 344.270 243.495 ;
        RECT 5.330 235.225 344.270 238.055 ;
        RECT 5.330 229.785 344.270 232.615 ;
        RECT 5.330 224.345 344.270 227.175 ;
        RECT 5.330 218.905 344.270 221.735 ;
        RECT 5.330 213.465 344.270 216.295 ;
        RECT 5.330 208.025 344.270 210.855 ;
        RECT 5.330 202.585 344.270 205.415 ;
        RECT 5.330 197.145 344.270 199.975 ;
        RECT 5.330 191.705 344.270 194.535 ;
        RECT 5.330 186.265 344.270 189.095 ;
        RECT 5.330 180.825 344.270 183.655 ;
        RECT 5.330 175.385 344.270 178.215 ;
        RECT 5.330 169.945 344.270 172.775 ;
        RECT 5.330 164.505 344.270 167.335 ;
        RECT 5.330 159.065 344.270 161.895 ;
        RECT 5.330 153.625 344.270 156.455 ;
        RECT 5.330 148.185 344.270 151.015 ;
        RECT 5.330 142.745 344.270 145.575 ;
        RECT 5.330 137.305 344.270 140.135 ;
        RECT 5.330 131.865 344.270 134.695 ;
        RECT 5.330 126.425 344.270 129.255 ;
        RECT 5.330 120.985 344.270 123.815 ;
        RECT 5.330 115.545 344.270 118.375 ;
        RECT 5.330 110.105 344.270 112.935 ;
        RECT 5.330 104.665 344.270 107.495 ;
        RECT 5.330 99.225 344.270 102.055 ;
        RECT 5.330 93.785 344.270 96.615 ;
        RECT 5.330 88.345 344.270 91.175 ;
        RECT 5.330 82.905 344.270 85.735 ;
        RECT 5.330 77.465 344.270 80.295 ;
        RECT 5.330 72.025 344.270 74.855 ;
        RECT 5.330 66.585 344.270 69.415 ;
        RECT 5.330 61.145 344.270 63.975 ;
        RECT 5.330 55.705 344.270 58.535 ;
        RECT 5.330 50.265 344.270 53.095 ;
        RECT 5.330 44.825 344.270 47.655 ;
        RECT 5.330 39.385 344.270 42.215 ;
        RECT 5.330 33.945 344.270 36.775 ;
        RECT 5.330 28.505 344.270 31.335 ;
        RECT 5.330 23.065 344.270 25.895 ;
        RECT 5.330 17.625 344.270 20.455 ;
        RECT 5.330 12.185 344.270 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 5.520 10.640 346.310 337.520 ;
      LAYER met2 ;
        RECT 7.000 10.695 346.280 337.465 ;
      LAYER met3 ;
        RECT 7.885 315.200 346.000 337.445 ;
        RECT 7.885 313.800 345.600 315.200 ;
        RECT 7.885 312.480 346.000 313.800 ;
        RECT 7.885 311.080 345.600 312.480 ;
        RECT 7.885 309.760 346.000 311.080 ;
        RECT 7.885 308.360 345.600 309.760 ;
        RECT 7.885 307.040 346.000 308.360 ;
        RECT 7.885 305.640 345.600 307.040 ;
        RECT 7.885 304.320 346.000 305.640 ;
        RECT 7.885 302.920 345.600 304.320 ;
        RECT 7.885 301.600 346.000 302.920 ;
        RECT 7.885 300.200 345.600 301.600 ;
        RECT 7.885 298.880 346.000 300.200 ;
        RECT 7.885 297.480 345.600 298.880 ;
        RECT 7.885 296.160 346.000 297.480 ;
        RECT 7.885 294.760 345.600 296.160 ;
        RECT 7.885 293.440 346.000 294.760 ;
        RECT 7.885 292.040 345.600 293.440 ;
        RECT 7.885 290.720 346.000 292.040 ;
        RECT 7.885 289.320 345.600 290.720 ;
        RECT 7.885 288.000 346.000 289.320 ;
        RECT 7.885 286.600 345.600 288.000 ;
        RECT 7.885 285.280 346.000 286.600 ;
        RECT 7.885 283.880 345.600 285.280 ;
        RECT 7.885 282.560 346.000 283.880 ;
        RECT 7.885 281.160 345.600 282.560 ;
        RECT 7.885 279.840 346.000 281.160 ;
        RECT 7.885 278.440 345.600 279.840 ;
        RECT 7.885 277.120 346.000 278.440 ;
        RECT 7.885 275.720 345.600 277.120 ;
        RECT 7.885 274.400 346.000 275.720 ;
        RECT 7.885 273.000 345.600 274.400 ;
        RECT 7.885 271.680 346.000 273.000 ;
        RECT 7.885 270.280 345.600 271.680 ;
        RECT 7.885 268.960 346.000 270.280 ;
        RECT 7.885 267.560 345.600 268.960 ;
        RECT 7.885 266.240 346.000 267.560 ;
        RECT 7.885 264.840 345.600 266.240 ;
        RECT 7.885 263.520 346.000 264.840 ;
        RECT 7.885 262.120 345.600 263.520 ;
        RECT 7.885 260.800 346.000 262.120 ;
        RECT 7.885 259.400 345.600 260.800 ;
        RECT 7.885 258.080 346.000 259.400 ;
        RECT 7.885 256.680 345.600 258.080 ;
        RECT 7.885 255.360 346.000 256.680 ;
        RECT 7.885 253.960 345.600 255.360 ;
        RECT 7.885 252.640 346.000 253.960 ;
        RECT 7.885 251.240 345.600 252.640 ;
        RECT 7.885 249.920 346.000 251.240 ;
        RECT 7.885 248.520 345.600 249.920 ;
        RECT 7.885 247.200 346.000 248.520 ;
        RECT 7.885 245.800 345.600 247.200 ;
        RECT 7.885 244.480 346.000 245.800 ;
        RECT 7.885 243.080 345.600 244.480 ;
        RECT 7.885 241.760 346.000 243.080 ;
        RECT 7.885 240.360 345.600 241.760 ;
        RECT 7.885 239.040 346.000 240.360 ;
        RECT 7.885 237.640 345.600 239.040 ;
        RECT 7.885 236.320 346.000 237.640 ;
        RECT 7.885 234.920 345.600 236.320 ;
        RECT 7.885 233.600 346.000 234.920 ;
        RECT 7.885 232.200 345.600 233.600 ;
        RECT 7.885 230.880 346.000 232.200 ;
        RECT 7.885 229.480 345.600 230.880 ;
        RECT 7.885 228.160 346.000 229.480 ;
        RECT 7.885 226.760 345.600 228.160 ;
        RECT 7.885 225.440 346.000 226.760 ;
        RECT 7.885 224.040 345.600 225.440 ;
        RECT 7.885 222.720 346.000 224.040 ;
        RECT 7.885 221.320 345.600 222.720 ;
        RECT 7.885 220.000 346.000 221.320 ;
        RECT 7.885 218.600 345.600 220.000 ;
        RECT 7.885 217.280 346.000 218.600 ;
        RECT 7.885 215.880 345.600 217.280 ;
        RECT 7.885 214.560 346.000 215.880 ;
        RECT 7.885 213.160 345.600 214.560 ;
        RECT 7.885 211.840 346.000 213.160 ;
        RECT 7.885 210.440 345.600 211.840 ;
        RECT 7.885 209.120 346.000 210.440 ;
        RECT 7.885 207.720 345.600 209.120 ;
        RECT 7.885 206.400 346.000 207.720 ;
        RECT 7.885 205.000 345.600 206.400 ;
        RECT 7.885 203.680 346.000 205.000 ;
        RECT 7.885 202.280 345.600 203.680 ;
        RECT 7.885 200.960 346.000 202.280 ;
        RECT 7.885 199.560 345.600 200.960 ;
        RECT 7.885 198.240 346.000 199.560 ;
        RECT 7.885 196.840 345.600 198.240 ;
        RECT 7.885 195.520 346.000 196.840 ;
        RECT 7.885 194.120 345.600 195.520 ;
        RECT 7.885 192.800 346.000 194.120 ;
        RECT 7.885 191.400 345.600 192.800 ;
        RECT 7.885 190.080 346.000 191.400 ;
        RECT 7.885 188.680 345.600 190.080 ;
        RECT 7.885 187.360 346.000 188.680 ;
        RECT 7.885 185.960 345.600 187.360 ;
        RECT 7.885 184.640 346.000 185.960 ;
        RECT 7.885 183.240 345.600 184.640 ;
        RECT 7.885 181.920 346.000 183.240 ;
        RECT 7.885 180.520 345.600 181.920 ;
        RECT 7.885 179.200 346.000 180.520 ;
        RECT 7.885 177.800 345.600 179.200 ;
        RECT 7.885 176.480 346.000 177.800 ;
        RECT 7.885 175.080 345.600 176.480 ;
        RECT 7.885 173.760 346.000 175.080 ;
        RECT 7.885 172.360 345.600 173.760 ;
        RECT 7.885 171.040 346.000 172.360 ;
        RECT 7.885 169.640 345.600 171.040 ;
        RECT 7.885 168.320 346.000 169.640 ;
        RECT 7.885 166.920 345.600 168.320 ;
        RECT 7.885 165.600 346.000 166.920 ;
        RECT 7.885 164.200 345.600 165.600 ;
        RECT 7.885 162.880 346.000 164.200 ;
        RECT 7.885 161.480 345.600 162.880 ;
        RECT 7.885 160.160 346.000 161.480 ;
        RECT 7.885 158.760 345.600 160.160 ;
        RECT 7.885 157.440 346.000 158.760 ;
        RECT 7.885 156.040 345.600 157.440 ;
        RECT 7.885 154.720 346.000 156.040 ;
        RECT 7.885 153.320 345.600 154.720 ;
        RECT 7.885 152.000 346.000 153.320 ;
        RECT 7.885 150.600 345.600 152.000 ;
        RECT 7.885 149.280 346.000 150.600 ;
        RECT 7.885 147.880 345.600 149.280 ;
        RECT 7.885 146.560 346.000 147.880 ;
        RECT 7.885 145.160 345.600 146.560 ;
        RECT 7.885 143.840 346.000 145.160 ;
        RECT 7.885 142.440 345.600 143.840 ;
        RECT 7.885 141.120 346.000 142.440 ;
        RECT 7.885 139.720 345.600 141.120 ;
        RECT 7.885 138.400 346.000 139.720 ;
        RECT 7.885 137.000 345.600 138.400 ;
        RECT 7.885 135.680 346.000 137.000 ;
        RECT 7.885 134.280 345.600 135.680 ;
        RECT 7.885 132.960 346.000 134.280 ;
        RECT 7.885 131.560 345.600 132.960 ;
        RECT 7.885 130.240 346.000 131.560 ;
        RECT 7.885 128.840 345.600 130.240 ;
        RECT 7.885 127.520 346.000 128.840 ;
        RECT 7.885 126.120 345.600 127.520 ;
        RECT 7.885 124.800 346.000 126.120 ;
        RECT 7.885 123.400 345.600 124.800 ;
        RECT 7.885 122.080 346.000 123.400 ;
        RECT 7.885 120.680 345.600 122.080 ;
        RECT 7.885 119.360 346.000 120.680 ;
        RECT 7.885 117.960 345.600 119.360 ;
        RECT 7.885 116.640 346.000 117.960 ;
        RECT 7.885 115.240 345.600 116.640 ;
        RECT 7.885 113.920 346.000 115.240 ;
        RECT 7.885 112.520 345.600 113.920 ;
        RECT 7.885 111.200 346.000 112.520 ;
        RECT 7.885 109.800 345.600 111.200 ;
        RECT 7.885 108.480 346.000 109.800 ;
        RECT 7.885 107.080 345.600 108.480 ;
        RECT 7.885 105.760 346.000 107.080 ;
        RECT 7.885 104.360 345.600 105.760 ;
        RECT 7.885 103.040 346.000 104.360 ;
        RECT 7.885 101.640 345.600 103.040 ;
        RECT 7.885 100.320 346.000 101.640 ;
        RECT 7.885 98.920 345.600 100.320 ;
        RECT 7.885 97.600 346.000 98.920 ;
        RECT 7.885 96.200 345.600 97.600 ;
        RECT 7.885 94.880 346.000 96.200 ;
        RECT 7.885 93.480 345.600 94.880 ;
        RECT 7.885 92.160 346.000 93.480 ;
        RECT 7.885 90.760 345.600 92.160 ;
        RECT 7.885 89.440 346.000 90.760 ;
        RECT 7.885 88.040 345.600 89.440 ;
        RECT 7.885 86.720 346.000 88.040 ;
        RECT 7.885 85.320 345.600 86.720 ;
        RECT 7.885 84.000 346.000 85.320 ;
        RECT 7.885 82.600 345.600 84.000 ;
        RECT 7.885 81.280 346.000 82.600 ;
        RECT 7.885 79.880 345.600 81.280 ;
        RECT 7.885 78.560 346.000 79.880 ;
        RECT 7.885 77.160 345.600 78.560 ;
        RECT 7.885 75.840 346.000 77.160 ;
        RECT 7.885 74.440 345.600 75.840 ;
        RECT 7.885 73.120 346.000 74.440 ;
        RECT 7.885 71.720 345.600 73.120 ;
        RECT 7.885 70.400 346.000 71.720 ;
        RECT 7.885 69.000 345.600 70.400 ;
        RECT 7.885 67.680 346.000 69.000 ;
        RECT 7.885 66.280 345.600 67.680 ;
        RECT 7.885 64.960 346.000 66.280 ;
        RECT 7.885 63.560 345.600 64.960 ;
        RECT 7.885 62.240 346.000 63.560 ;
        RECT 7.885 60.840 345.600 62.240 ;
        RECT 7.885 59.520 346.000 60.840 ;
        RECT 7.885 58.120 345.600 59.520 ;
        RECT 7.885 56.800 346.000 58.120 ;
        RECT 7.885 55.400 345.600 56.800 ;
        RECT 7.885 54.080 346.000 55.400 ;
        RECT 7.885 52.680 345.600 54.080 ;
        RECT 7.885 51.360 346.000 52.680 ;
        RECT 7.885 49.960 345.600 51.360 ;
        RECT 7.885 48.640 346.000 49.960 ;
        RECT 7.885 47.240 345.600 48.640 ;
        RECT 7.885 45.920 346.000 47.240 ;
        RECT 7.885 44.520 345.600 45.920 ;
        RECT 7.885 43.200 346.000 44.520 ;
        RECT 7.885 41.800 345.600 43.200 ;
        RECT 7.885 40.480 346.000 41.800 ;
        RECT 7.885 39.080 345.600 40.480 ;
        RECT 7.885 37.760 346.000 39.080 ;
        RECT 7.885 36.360 345.600 37.760 ;
        RECT 7.885 35.040 346.000 36.360 ;
        RECT 7.885 33.640 345.600 35.040 ;
        RECT 7.885 10.715 346.000 33.640 ;
      LAYER met4 ;
        RECT 67.455 19.895 97.440 331.665 ;
        RECT 99.840 19.895 174.240 331.665 ;
        RECT 176.640 19.895 251.040 331.665 ;
        RECT 253.440 19.895 327.840 331.665 ;
        RECT 330.240 19.895 337.345 331.665 ;
      LAYER met5 ;
        RECT 81.540 65.500 318.660 254.100 ;
  END
END alu
END LIBRARY

