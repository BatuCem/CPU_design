VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO datapath
  CLASS BLOCK ;
  FOREIGN datapath ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN ALUASrcSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.840 400.000 143.440 ;
    END
  END ALUASrcSel
  PIN ALUBSrcSel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END ALUBSrcSel[0]
  PIN ALUBSrcSel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END ALUBSrcSel[1]
  PIN AluResult[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END AluResult[0]
  PIN AluResult[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END AluResult[10]
  PIN AluResult[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END AluResult[11]
  PIN AluResult[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END AluResult[12]
  PIN AluResult[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END AluResult[13]
  PIN AluResult[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END AluResult[14]
  PIN AluResult[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END AluResult[15]
  PIN AluResult[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END AluResult[16]
  PIN AluResult[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END AluResult[17]
  PIN AluResult[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END AluResult[18]
  PIN AluResult[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END AluResult[19]
  PIN AluResult[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END AluResult[1]
  PIN AluResult[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END AluResult[20]
  PIN AluResult[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END AluResult[21]
  PIN AluResult[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END AluResult[22]
  PIN AluResult[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END AluResult[23]
  PIN AluResult[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END AluResult[24]
  PIN AluResult[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END AluResult[25]
  PIN AluResult[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END AluResult[26]
  PIN AluResult[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END AluResult[27]
  PIN AluResult[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END AluResult[28]
  PIN AluResult[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END AluResult[29]
  PIN AluResult[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END AluResult[2]
  PIN AluResult[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END AluResult[30]
  PIN AluResult[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END AluResult[31]
  PIN AluResult[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END AluResult[3]
  PIN AluResult[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END AluResult[4]
  PIN AluResult[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END AluResult[5]
  PIN AluResult[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END AluResult[6]
  PIN AluResult[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END AluResult[7]
  PIN AluResult[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END AluResult[8]
  PIN AluResult[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END AluResult[9]
  PIN IRWriteEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 153.720 400.000 154.320 ;
    END
  END IRWriteEn
  PIN IorDSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.000 400.000 151.600 ;
    END
  END IorDSel
  PIN MemtoRegSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 140.120 400.000 140.720 ;
    END
  END MemtoRegSel
  PIN PCEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END PCEn
  PIN PCSrcSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 148.280 400.000 148.880 ;
    END
  END PCSrcSel
  PIN RegDstSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 145.560 400.000 146.160 ;
    END
  END RegDstSel
  PIN SrcA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END SrcA[0]
  PIN SrcA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END SrcA[10]
  PIN SrcA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END SrcA[11]
  PIN SrcA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END SrcA[12]
  PIN SrcA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END SrcA[13]
  PIN SrcA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END SrcA[14]
  PIN SrcA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END SrcA[15]
  PIN SrcA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END SrcA[16]
  PIN SrcA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END SrcA[17]
  PIN SrcA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END SrcA[18]
  PIN SrcA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END SrcA[19]
  PIN SrcA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END SrcA[1]
  PIN SrcA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END SrcA[20]
  PIN SrcA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END SrcA[21]
  PIN SrcA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END SrcA[22]
  PIN SrcA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END SrcA[23]
  PIN SrcA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END SrcA[24]
  PIN SrcA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END SrcA[25]
  PIN SrcA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END SrcA[26]
  PIN SrcA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END SrcA[27]
  PIN SrcA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END SrcA[28]
  PIN SrcA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END SrcA[29]
  PIN SrcA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END SrcA[2]
  PIN SrcA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END SrcA[30]
  PIN SrcA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END SrcA[31]
  PIN SrcA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END SrcA[3]
  PIN SrcA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END SrcA[4]
  PIN SrcA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END SrcA[5]
  PIN SrcA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END SrcA[6]
  PIN SrcA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END SrcA[7]
  PIN SrcA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END SrcA[8]
  PIN SrcA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END SrcA[9]
  PIN SrcB[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END SrcB[0]
  PIN SrcB[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END SrcB[10]
  PIN SrcB[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END SrcB[11]
  PIN SrcB[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END SrcB[12]
  PIN SrcB[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END SrcB[13]
  PIN SrcB[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END SrcB[14]
  PIN SrcB[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END SrcB[15]
  PIN SrcB[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END SrcB[16]
  PIN SrcB[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END SrcB[17]
  PIN SrcB[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END SrcB[18]
  PIN SrcB[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END SrcB[19]
  PIN SrcB[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END SrcB[1]
  PIN SrcB[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END SrcB[20]
  PIN SrcB[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END SrcB[21]
  PIN SrcB[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END SrcB[22]
  PIN SrcB[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END SrcB[23]
  PIN SrcB[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END SrcB[24]
  PIN SrcB[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END SrcB[25]
  PIN SrcB[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END SrcB[26]
  PIN SrcB[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END SrcB[27]
  PIN SrcB[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END SrcB[28]
  PIN SrcB[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END SrcB[29]
  PIN SrcB[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END SrcB[2]
  PIN SrcB[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END SrcB[30]
  PIN SrcB[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END SrcB[31]
  PIN SrcB[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END SrcB[3]
  PIN SrcB[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END SrcB[4]
  PIN SrcB[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END SrcB[5]
  PIN SrcB[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END SrcB[6]
  PIN SrcB[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END SrcB[7]
  PIN SrcB[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END SrcB[8]
  PIN SrcB[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END SrcB[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END VPWR
  PIN addr_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 98.990 396.000 99.270 400.000 ;
    END
  END addr_mem[0]
  PIN addr_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 126.590 396.000 126.870 400.000 ;
    END
  END addr_mem[10]
  PIN addr_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 129.350 396.000 129.630 400.000 ;
    END
  END addr_mem[11]
  PIN addr_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 396.000 132.390 400.000 ;
    END
  END addr_mem[12]
  PIN addr_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 134.870 396.000 135.150 400.000 ;
    END
  END addr_mem[13]
  PIN addr_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 137.630 396.000 137.910 400.000 ;
    END
  END addr_mem[14]
  PIN addr_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 140.390 396.000 140.670 400.000 ;
    END
  END addr_mem[15]
  PIN addr_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 143.150 396.000 143.430 400.000 ;
    END
  END addr_mem[16]
  PIN addr_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 145.910 396.000 146.190 400.000 ;
    END
  END addr_mem[17]
  PIN addr_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.670 396.000 148.950 400.000 ;
    END
  END addr_mem[18]
  PIN addr_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 396.000 151.710 400.000 ;
    END
  END addr_mem[19]
  PIN addr_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 101.750 396.000 102.030 400.000 ;
    END
  END addr_mem[1]
  PIN addr_mem[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 154.190 396.000 154.470 400.000 ;
    END
  END addr_mem[20]
  PIN addr_mem[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 156.950 396.000 157.230 400.000 ;
    END
  END addr_mem[21]
  PIN addr_mem[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 159.710 396.000 159.990 400.000 ;
    END
  END addr_mem[22]
  PIN addr_mem[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.470 396.000 162.750 400.000 ;
    END
  END addr_mem[23]
  PIN addr_mem[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 165.230 396.000 165.510 400.000 ;
    END
  END addr_mem[24]
  PIN addr_mem[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.990 396.000 168.270 400.000 ;
    END
  END addr_mem[25]
  PIN addr_mem[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 170.750 396.000 171.030 400.000 ;
    END
  END addr_mem[26]
  PIN addr_mem[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 173.510 396.000 173.790 400.000 ;
    END
  END addr_mem[27]
  PIN addr_mem[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 176.270 396.000 176.550 400.000 ;
    END
  END addr_mem[28]
  PIN addr_mem[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 179.030 396.000 179.310 400.000 ;
    END
  END addr_mem[29]
  PIN addr_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 104.510 396.000 104.790 400.000 ;
    END
  END addr_mem[2]
  PIN addr_mem[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 181.790 396.000 182.070 400.000 ;
    END
  END addr_mem[30]
  PIN addr_mem[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 184.550 396.000 184.830 400.000 ;
    END
  END addr_mem[31]
  PIN addr_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 396.000 107.550 400.000 ;
    END
  END addr_mem[3]
  PIN addr_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 110.030 396.000 110.310 400.000 ;
    END
  END addr_mem[4]
  PIN addr_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 112.790 396.000 113.070 400.000 ;
    END
  END addr_mem[5]
  PIN addr_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 115.550 396.000 115.830 400.000 ;
    END
  END addr_mem[6]
  PIN addr_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 118.310 396.000 118.590 400.000 ;
    END
  END addr_mem[7]
  PIN addr_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 121.070 396.000 121.350 400.000 ;
    END
  END addr_mem[8]
  PIN addr_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 123.830 396.000 124.110 400.000 ;
    END
  END addr_mem[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END clk
  PIN instruction[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 275.630 396.000 275.910 400.000 ;
    END
  END instruction[0]
  PIN instruction[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 303.230 396.000 303.510 400.000 ;
    END
  END instruction[10]
  PIN instruction[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 305.990 396.000 306.270 400.000 ;
    END
  END instruction[11]
  PIN instruction[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 308.750 396.000 309.030 400.000 ;
    END
  END instruction[12]
  PIN instruction[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 311.510 396.000 311.790 400.000 ;
    END
  END instruction[13]
  PIN instruction[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 314.270 396.000 314.550 400.000 ;
    END
  END instruction[14]
  PIN instruction[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 317.030 396.000 317.310 400.000 ;
    END
  END instruction[15]
  PIN instruction[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 319.790 396.000 320.070 400.000 ;
    END
  END instruction[16]
  PIN instruction[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 322.550 396.000 322.830 400.000 ;
    END
  END instruction[17]
  PIN instruction[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 396.000 325.590 400.000 ;
    END
  END instruction[18]
  PIN instruction[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 328.070 396.000 328.350 400.000 ;
    END
  END instruction[19]
  PIN instruction[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 278.390 396.000 278.670 400.000 ;
    END
  END instruction[1]
  PIN instruction[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 330.830 396.000 331.110 400.000 ;
    END
  END instruction[20]
  PIN instruction[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 333.590 396.000 333.870 400.000 ;
    END
  END instruction[21]
  PIN instruction[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 336.350 396.000 336.630 400.000 ;
    END
  END instruction[22]
  PIN instruction[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 339.110 396.000 339.390 400.000 ;
    END
  END instruction[23]
  PIN instruction[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 341.870 396.000 342.150 400.000 ;
    END
  END instruction[24]
  PIN instruction[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 344.630 396.000 344.910 400.000 ;
    END
  END instruction[25]
  PIN instruction[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 347.390 396.000 347.670 400.000 ;
    END
  END instruction[26]
  PIN instruction[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 350.150 396.000 350.430 400.000 ;
    END
  END instruction[27]
  PIN instruction[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 352.910 396.000 353.190 400.000 ;
    END
  END instruction[28]
  PIN instruction[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 355.670 396.000 355.950 400.000 ;
    END
  END instruction[29]
  PIN instruction[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 281.150 396.000 281.430 400.000 ;
    END
  END instruction[2]
  PIN instruction[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 358.430 396.000 358.710 400.000 ;
    END
  END instruction[30]
  PIN instruction[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 361.190 396.000 361.470 400.000 ;
    END
  END instruction[31]
  PIN instruction[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 283.910 396.000 284.190 400.000 ;
    END
  END instruction[3]
  PIN instruction[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 396.000 286.950 400.000 ;
    END
  END instruction[4]
  PIN instruction[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 289.430 396.000 289.710 400.000 ;
    END
  END instruction[5]
  PIN instruction[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 292.190 396.000 292.470 400.000 ;
    END
  END instruction[6]
  PIN instruction[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 294.950 396.000 295.230 400.000 ;
    END
  END instruction[7]
  PIN instruction[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 297.710 396.000 297.990 400.000 ;
    END
  END instruction[8]
  PIN instruction[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 300.470 396.000 300.750 400.000 ;
    END
  END instruction[9]
  PIN mem_Wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 10.670 396.000 10.950 400.000 ;
    END
  END mem_Wdata[0]
  PIN mem_Wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.270 396.000 38.550 400.000 ;
    END
  END mem_Wdata[10]
  PIN mem_Wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.030 396.000 41.310 400.000 ;
    END
  END mem_Wdata[11]
  PIN mem_Wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 43.790 396.000 44.070 400.000 ;
    END
  END mem_Wdata[12]
  PIN mem_Wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 46.550 396.000 46.830 400.000 ;
    END
  END mem_Wdata[13]
  PIN mem_Wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 49.310 396.000 49.590 400.000 ;
    END
  END mem_Wdata[14]
  PIN mem_Wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.070 396.000 52.350 400.000 ;
    END
  END mem_Wdata[15]
  PIN mem_Wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 396.000 55.110 400.000 ;
    END
  END mem_Wdata[16]
  PIN mem_Wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 57.590 396.000 57.870 400.000 ;
    END
  END mem_Wdata[17]
  PIN mem_Wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 60.350 396.000 60.630 400.000 ;
    END
  END mem_Wdata[18]
  PIN mem_Wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 63.110 396.000 63.390 400.000 ;
    END
  END mem_Wdata[19]
  PIN mem_Wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 13.430 396.000 13.710 400.000 ;
    END
  END mem_Wdata[1]
  PIN mem_Wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.870 396.000 66.150 400.000 ;
    END
  END mem_Wdata[20]
  PIN mem_Wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 68.630 396.000 68.910 400.000 ;
    END
  END mem_Wdata[21]
  PIN mem_Wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 71.390 396.000 71.670 400.000 ;
    END
  END mem_Wdata[22]
  PIN mem_Wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 396.000 74.430 400.000 ;
    END
  END mem_Wdata[23]
  PIN mem_Wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 76.910 396.000 77.190 400.000 ;
    END
  END mem_Wdata[24]
  PIN mem_Wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 79.670 396.000 79.950 400.000 ;
    END
  END mem_Wdata[25]
  PIN mem_Wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.430 396.000 82.710 400.000 ;
    END
  END mem_Wdata[26]
  PIN mem_Wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 85.190 396.000 85.470 400.000 ;
    END
  END mem_Wdata[27]
  PIN mem_Wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.950 396.000 88.230 400.000 ;
    END
  END mem_Wdata[28]
  PIN mem_Wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.710 396.000 90.990 400.000 ;
    END
  END mem_Wdata[29]
  PIN mem_Wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 396.000 16.470 400.000 ;
    END
  END mem_Wdata[2]
  PIN mem_Wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 396.000 93.750 400.000 ;
    END
  END mem_Wdata[30]
  PIN mem_Wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.230 396.000 96.510 400.000 ;
    END
  END mem_Wdata[31]
  PIN mem_Wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 18.950 396.000 19.230 400.000 ;
    END
  END mem_Wdata[3]
  PIN mem_Wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 21.710 396.000 21.990 400.000 ;
    END
  END mem_Wdata[4]
  PIN mem_Wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 24.470 396.000 24.750 400.000 ;
    END
  END mem_Wdata[5]
  PIN mem_Wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 27.230 396.000 27.510 400.000 ;
    END
  END mem_Wdata[6]
  PIN mem_Wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.990 396.000 30.270 400.000 ;
    END
  END mem_Wdata[7]
  PIN mem_Wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.750 396.000 33.030 400.000 ;
    END
  END mem_Wdata[8]
  PIN mem_Wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 396.000 35.790 400.000 ;
    END
  END mem_Wdata[9]
  PIN override_memread
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END override_memread
  PIN override_memwrite
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END override_memwrite
  PIN override_rwaddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END override_rwaddr[0]
  PIN override_rwaddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END override_rwaddr[10]
  PIN override_rwaddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END override_rwaddr[11]
  PIN override_rwaddr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END override_rwaddr[12]
  PIN override_rwaddr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END override_rwaddr[13]
  PIN override_rwaddr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END override_rwaddr[14]
  PIN override_rwaddr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END override_rwaddr[15]
  PIN override_rwaddr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END override_rwaddr[16]
  PIN override_rwaddr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END override_rwaddr[17]
  PIN override_rwaddr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END override_rwaddr[18]
  PIN override_rwaddr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END override_rwaddr[19]
  PIN override_rwaddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END override_rwaddr[1]
  PIN override_rwaddr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END override_rwaddr[20]
  PIN override_rwaddr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END override_rwaddr[21]
  PIN override_rwaddr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END override_rwaddr[22]
  PIN override_rwaddr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END override_rwaddr[23]
  PIN override_rwaddr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END override_rwaddr[24]
  PIN override_rwaddr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END override_rwaddr[25]
  PIN override_rwaddr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END override_rwaddr[26]
  PIN override_rwaddr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END override_rwaddr[27]
  PIN override_rwaddr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END override_rwaddr[28]
  PIN override_rwaddr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END override_rwaddr[29]
  PIN override_rwaddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END override_rwaddr[2]
  PIN override_rwaddr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END override_rwaddr[30]
  PIN override_rwaddr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END override_rwaddr[31]
  PIN override_rwaddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END override_rwaddr[3]
  PIN override_rwaddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END override_rwaddr[4]
  PIN override_rwaddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END override_rwaddr[5]
  PIN override_rwaddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END override_rwaddr[6]
  PIN override_rwaddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END override_rwaddr[7]
  PIN override_rwaddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END override_rwaddr[8]
  PIN override_rwaddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END override_rwaddr[9]
  PIN override_rwdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END override_rwdata[0]
  PIN override_rwdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END override_rwdata[10]
  PIN override_rwdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END override_rwdata[11]
  PIN override_rwdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END override_rwdata[12]
  PIN override_rwdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END override_rwdata[13]
  PIN override_rwdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END override_rwdata[14]
  PIN override_rwdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END override_rwdata[15]
  PIN override_rwdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END override_rwdata[16]
  PIN override_rwdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END override_rwdata[17]
  PIN override_rwdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END override_rwdata[18]
  PIN override_rwdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END override_rwdata[19]
  PIN override_rwdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END override_rwdata[1]
  PIN override_rwdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END override_rwdata[20]
  PIN override_rwdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END override_rwdata[21]
  PIN override_rwdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END override_rwdata[22]
  PIN override_rwdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END override_rwdata[23]
  PIN override_rwdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END override_rwdata[24]
  PIN override_rwdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END override_rwdata[25]
  PIN override_rwdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END override_rwdata[26]
  PIN override_rwdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END override_rwdata[27]
  PIN override_rwdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END override_rwdata[28]
  PIN override_rwdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END override_rwdata[29]
  PIN override_rwdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END override_rwdata[2]
  PIN override_rwdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END override_rwdata[30]
  PIN override_rwdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END override_rwdata[31]
  PIN override_rwdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END override_rwdata[3]
  PIN override_rwdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END override_rwdata[4]
  PIN override_rwdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END override_rwdata[5]
  PIN override_rwdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END override_rwdata[6]
  PIN override_rwdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END override_rwdata[7]
  PIN override_rwdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END override_rwdata[8]
  PIN override_rwdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END override_rwdata[9]
  PIN regA2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 363.950 396.000 364.230 400.000 ;
    END
  END regA2[0]
  PIN regA2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 366.710 396.000 366.990 400.000 ;
    END
  END regA2[1]
  PIN regA2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 369.470 396.000 369.750 400.000 ;
    END
  END regA2[2]
  PIN regA2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 372.230 396.000 372.510 400.000 ;
    END
  END regA2[3]
  PIN regA2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 374.990 396.000 375.270 400.000 ;
    END
  END regA2[4]
  PIN regA3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 377.750 396.000 378.030 400.000 ;
    END
  END regA3[0]
  PIN regA3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 380.510 396.000 380.790 400.000 ;
    END
  END regA3[1]
  PIN regA3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 396.000 383.550 400.000 ;
    END
  END regA3[2]
  PIN regA3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 386.030 396.000 386.310 400.000 ;
    END
  END regA3[3]
  PIN regA3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 388.790 396.000 389.070 400.000 ;
    END
  END regA3[4]
  PIN reg_instr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 53.080 400.000 53.680 ;
    END
  END reg_instr[0]
  PIN reg_instr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 80.280 400.000 80.880 ;
    END
  END reg_instr[10]
  PIN reg_instr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 83.000 400.000 83.600 ;
    END
  END reg_instr[11]
  PIN reg_instr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.720 400.000 86.320 ;
    END
  END reg_instr[12]
  PIN reg_instr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 88.440 400.000 89.040 ;
    END
  END reg_instr[13]
  PIN reg_instr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.160 400.000 91.760 ;
    END
  END reg_instr[14]
  PIN reg_instr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 93.880 400.000 94.480 ;
    END
  END reg_instr[15]
  PIN reg_instr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 96.600 400.000 97.200 ;
    END
  END reg_instr[16]
  PIN reg_instr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 99.320 400.000 99.920 ;
    END
  END reg_instr[17]
  PIN reg_instr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.040 400.000 102.640 ;
    END
  END reg_instr[18]
  PIN reg_instr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.760 400.000 105.360 ;
    END
  END reg_instr[19]
  PIN reg_instr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 55.800 400.000 56.400 ;
    END
  END reg_instr[1]
  PIN reg_instr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 107.480 400.000 108.080 ;
    END
  END reg_instr[20]
  PIN reg_instr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 110.200 400.000 110.800 ;
    END
  END reg_instr[21]
  PIN reg_instr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.920 400.000 113.520 ;
    END
  END reg_instr[22]
  PIN reg_instr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 115.640 400.000 116.240 ;
    END
  END reg_instr[23]
  PIN reg_instr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 118.360 400.000 118.960 ;
    END
  END reg_instr[24]
  PIN reg_instr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 121.080 400.000 121.680 ;
    END
  END reg_instr[25]
  PIN reg_instr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.800 400.000 124.400 ;
    END
  END reg_instr[26]
  PIN reg_instr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 126.520 400.000 127.120 ;
    END
  END reg_instr[27]
  PIN reg_instr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.240 400.000 129.840 ;
    END
  END reg_instr[28]
  PIN reg_instr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 131.960 400.000 132.560 ;
    END
  END reg_instr[29]
  PIN reg_instr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 58.520 400.000 59.120 ;
    END
  END reg_instr[2]
  PIN reg_instr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 134.680 400.000 135.280 ;
    END
  END reg_instr[30]
  PIN reg_instr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 137.400 400.000 138.000 ;
    END
  END reg_instr[31]
  PIN reg_instr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.240 400.000 61.840 ;
    END
  END reg_instr[3]
  PIN reg_instr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 63.960 400.000 64.560 ;
    END
  END reg_instr[4]
  PIN reg_instr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 66.680 400.000 67.280 ;
    END
  END reg_instr[5]
  PIN reg_instr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 69.400 400.000 70.000 ;
    END
  END reg_instr[6]
  PIN reg_instr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.120 400.000 72.720 ;
    END
  END reg_instr[7]
  PIN reg_instr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.840 400.000 75.440 ;
    END
  END reg_instr[8]
  PIN reg_instr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 77.560 400.000 78.160 ;
    END
  END reg_instr[9]
  PIN reg_writeaddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.240 400.000 333.840 ;
    END
  END reg_writeaddr[0]
  PIN reg_writeaddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 335.960 400.000 336.560 ;
    END
  END reg_writeaddr[1]
  PIN reg_writeaddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 338.680 400.000 339.280 ;
    END
  END reg_writeaddr[2]
  PIN reg_writeaddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 341.400 400.000 342.000 ;
    END
  END reg_writeaddr[3]
  PIN reg_writeaddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 396.000 344.120 400.000 344.720 ;
    END
  END reg_writeaddr[4]
  PIN reg_writedata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 187.310 396.000 187.590 400.000 ;
    END
  END reg_writedata[0]
  PIN reg_writedata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 214.910 396.000 215.190 400.000 ;
    END
  END reg_writedata[10]
  PIN reg_writedata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 217.670 396.000 217.950 400.000 ;
    END
  END reg_writedata[11]
  PIN reg_writedata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 220.430 396.000 220.710 400.000 ;
    END
  END reg_writedata[12]
  PIN reg_writedata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 223.190 396.000 223.470 400.000 ;
    END
  END reg_writedata[13]
  PIN reg_writedata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 225.950 396.000 226.230 400.000 ;
    END
  END reg_writedata[14]
  PIN reg_writedata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 228.710 396.000 228.990 400.000 ;
    END
  END reg_writedata[15]
  PIN reg_writedata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 231.470 396.000 231.750 400.000 ;
    END
  END reg_writedata[16]
  PIN reg_writedata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 234.230 396.000 234.510 400.000 ;
    END
  END reg_writedata[17]
  PIN reg_writedata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 236.990 396.000 237.270 400.000 ;
    END
  END reg_writedata[18]
  PIN reg_writedata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 239.750 396.000 240.030 400.000 ;
    END
  END reg_writedata[19]
  PIN reg_writedata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.070 396.000 190.350 400.000 ;
    END
  END reg_writedata[1]
  PIN reg_writedata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 242.510 396.000 242.790 400.000 ;
    END
  END reg_writedata[20]
  PIN reg_writedata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 245.270 396.000 245.550 400.000 ;
    END
  END reg_writedata[21]
  PIN reg_writedata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 248.030 396.000 248.310 400.000 ;
    END
  END reg_writedata[22]
  PIN reg_writedata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 250.790 396.000 251.070 400.000 ;
    END
  END reg_writedata[23]
  PIN reg_writedata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 253.550 396.000 253.830 400.000 ;
    END
  END reg_writedata[24]
  PIN reg_writedata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 256.310 396.000 256.590 400.000 ;
    END
  END reg_writedata[25]
  PIN reg_writedata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 259.070 396.000 259.350 400.000 ;
    END
  END reg_writedata[26]
  PIN reg_writedata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 261.830 396.000 262.110 400.000 ;
    END
  END reg_writedata[27]
  PIN reg_writedata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 264.590 396.000 264.870 400.000 ;
    END
  END reg_writedata[28]
  PIN reg_writedata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 267.350 396.000 267.630 400.000 ;
    END
  END reg_writedata[29]
  PIN reg_writedata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 192.830 396.000 193.110 400.000 ;
    END
  END reg_writedata[2]
  PIN reg_writedata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.110 396.000 270.390 400.000 ;
    END
  END reg_writedata[30]
  PIN reg_writedata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 272.870 396.000 273.150 400.000 ;
    END
  END reg_writedata[31]
  PIN reg_writedata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 195.590 396.000 195.870 400.000 ;
    END
  END reg_writedata[3]
  PIN reg_writedata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 198.350 396.000 198.630 400.000 ;
    END
  END reg_writedata[4]
  PIN reg_writedata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 201.110 396.000 201.390 400.000 ;
    END
  END reg_writedata[5]
  PIN reg_writedata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 203.870 396.000 204.150 400.000 ;
    END
  END reg_writedata[6]
  PIN reg_writedata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 206.630 396.000 206.910 400.000 ;
    END
  END reg_writedata[7]
  PIN reg_writedata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 209.390 396.000 209.670 400.000 ;
    END
  END reg_writedata[8]
  PIN reg_writedata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 212.150 396.000 212.430 400.000 ;
    END
  END reg_writedata[9]
  PIN regfile_readA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.160 400.000 159.760 ;
    END
  END regfile_readA[0]
  PIN regfile_readA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 186.360 400.000 186.960 ;
    END
  END regfile_readA[10]
  PIN regfile_readA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 189.080 400.000 189.680 ;
    END
  END regfile_readA[11]
  PIN regfile_readA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 191.800 400.000 192.400 ;
    END
  END regfile_readA[12]
  PIN regfile_readA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 194.520 400.000 195.120 ;
    END
  END regfile_readA[13]
  PIN regfile_readA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END regfile_readA[14]
  PIN regfile_readA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 199.960 400.000 200.560 ;
    END
  END regfile_readA[15]
  PIN regfile_readA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.680 400.000 203.280 ;
    END
  END regfile_readA[16]
  PIN regfile_readA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 205.400 400.000 206.000 ;
    END
  END regfile_readA[17]
  PIN regfile_readA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 208.120 400.000 208.720 ;
    END
  END regfile_readA[18]
  PIN regfile_readA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.840 400.000 211.440 ;
    END
  END regfile_readA[19]
  PIN regfile_readA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 161.880 400.000 162.480 ;
    END
  END regfile_readA[1]
  PIN regfile_readA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 213.560 400.000 214.160 ;
    END
  END regfile_readA[20]
  PIN regfile_readA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.280 400.000 216.880 ;
    END
  END regfile_readA[21]
  PIN regfile_readA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 219.000 400.000 219.600 ;
    END
  END regfile_readA[22]
  PIN regfile_readA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.720 400.000 222.320 ;
    END
  END regfile_readA[23]
  PIN regfile_readA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 224.440 400.000 225.040 ;
    END
  END regfile_readA[24]
  PIN regfile_readA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.160 400.000 227.760 ;
    END
  END regfile_readA[25]
  PIN regfile_readA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.880 400.000 230.480 ;
    END
  END regfile_readA[26]
  PIN regfile_readA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 232.600 400.000 233.200 ;
    END
  END regfile_readA[27]
  PIN regfile_readA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 235.320 400.000 235.920 ;
    END
  END regfile_readA[28]
  PIN regfile_readA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 400.000 238.640 ;
    END
  END regfile_readA[29]
  PIN regfile_readA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 164.600 400.000 165.200 ;
    END
  END regfile_readA[2]
  PIN regfile_readA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 240.760 400.000 241.360 ;
    END
  END regfile_readA[30]
  PIN regfile_readA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 243.480 400.000 244.080 ;
    END
  END regfile_readA[31]
  PIN regfile_readA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 167.320 400.000 167.920 ;
    END
  END regfile_readA[3]
  PIN regfile_readA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 400.000 170.640 ;
    END
  END regfile_readA[4]
  PIN regfile_readA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.760 400.000 173.360 ;
    END
  END regfile_readA[5]
  PIN regfile_readA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 175.480 400.000 176.080 ;
    END
  END regfile_readA[6]
  PIN regfile_readA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 178.200 400.000 178.800 ;
    END
  END regfile_readA[7]
  PIN regfile_readA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.920 400.000 181.520 ;
    END
  END regfile_readA[8]
  PIN regfile_readA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 183.640 400.000 184.240 ;
    END
  END regfile_readA[9]
  PIN regfile_readB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 246.200 400.000 246.800 ;
    END
  END regfile_readB[0]
  PIN regfile_readB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 273.400 400.000 274.000 ;
    END
  END regfile_readB[10]
  PIN regfile_readB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 276.120 400.000 276.720 ;
    END
  END regfile_readB[11]
  PIN regfile_readB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.840 400.000 279.440 ;
    END
  END regfile_readB[12]
  PIN regfile_readB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 281.560 400.000 282.160 ;
    END
  END regfile_readB[13]
  PIN regfile_readB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 284.280 400.000 284.880 ;
    END
  END regfile_readB[14]
  PIN regfile_readB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 287.000 400.000 287.600 ;
    END
  END regfile_readB[15]
  PIN regfile_readB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.720 400.000 290.320 ;
    END
  END regfile_readB[16]
  PIN regfile_readB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 292.440 400.000 293.040 ;
    END
  END regfile_readB[17]
  PIN regfile_readB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.160 400.000 295.760 ;
    END
  END regfile_readB[18]
  PIN regfile_readB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 297.880 400.000 298.480 ;
    END
  END regfile_readB[19]
  PIN regfile_readB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.920 400.000 249.520 ;
    END
  END regfile_readB[1]
  PIN regfile_readB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 300.600 400.000 301.200 ;
    END
  END regfile_readB[20]
  PIN regfile_readB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 303.320 400.000 303.920 ;
    END
  END regfile_readB[21]
  PIN regfile_readB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 400.000 306.640 ;
    END
  END regfile_readB[22]
  PIN regfile_readB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 308.760 400.000 309.360 ;
    END
  END regfile_readB[23]
  PIN regfile_readB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 311.480 400.000 312.080 ;
    END
  END regfile_readB[24]
  PIN regfile_readB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 314.200 400.000 314.800 ;
    END
  END regfile_readB[25]
  PIN regfile_readB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 316.920 400.000 317.520 ;
    END
  END regfile_readB[26]
  PIN regfile_readB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 319.640 400.000 320.240 ;
    END
  END regfile_readB[27]
  PIN regfile_readB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 322.360 400.000 322.960 ;
    END
  END regfile_readB[28]
  PIN regfile_readB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 325.080 400.000 325.680 ;
    END
  END regfile_readB[29]
  PIN regfile_readB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 251.640 400.000 252.240 ;
    END
  END regfile_readB[2]
  PIN regfile_readB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 327.800 400.000 328.400 ;
    END
  END regfile_readB[30]
  PIN regfile_readB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 330.520 400.000 331.120 ;
    END
  END regfile_readB[31]
  PIN regfile_readB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 254.360 400.000 254.960 ;
    END
  END regfile_readB[3]
  PIN regfile_readB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 257.080 400.000 257.680 ;
    END
  END regfile_readB[4]
  PIN regfile_readB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 259.800 400.000 260.400 ;
    END
  END regfile_readB[5]
  PIN regfile_readB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 262.520 400.000 263.120 ;
    END
  END regfile_readB[6]
  PIN regfile_readB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.240 400.000 265.840 ;
    END
  END regfile_readB[7]
  PIN regfile_readB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 267.960 400.000 268.560 ;
    END
  END regfile_readB[8]
  PIN regfile_readB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 270.680 400.000 271.280 ;
    END
  END regfile_readB[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 389.045 ;
      LAYER met1 ;
        RECT 4.670 10.640 395.530 391.300 ;
      LAYER met2 ;
        RECT 4.690 395.720 10.390 396.170 ;
        RECT 11.230 395.720 13.150 396.170 ;
        RECT 13.990 395.720 15.910 396.170 ;
        RECT 16.750 395.720 18.670 396.170 ;
        RECT 19.510 395.720 21.430 396.170 ;
        RECT 22.270 395.720 24.190 396.170 ;
        RECT 25.030 395.720 26.950 396.170 ;
        RECT 27.790 395.720 29.710 396.170 ;
        RECT 30.550 395.720 32.470 396.170 ;
        RECT 33.310 395.720 35.230 396.170 ;
        RECT 36.070 395.720 37.990 396.170 ;
        RECT 38.830 395.720 40.750 396.170 ;
        RECT 41.590 395.720 43.510 396.170 ;
        RECT 44.350 395.720 46.270 396.170 ;
        RECT 47.110 395.720 49.030 396.170 ;
        RECT 49.870 395.720 51.790 396.170 ;
        RECT 52.630 395.720 54.550 396.170 ;
        RECT 55.390 395.720 57.310 396.170 ;
        RECT 58.150 395.720 60.070 396.170 ;
        RECT 60.910 395.720 62.830 396.170 ;
        RECT 63.670 395.720 65.590 396.170 ;
        RECT 66.430 395.720 68.350 396.170 ;
        RECT 69.190 395.720 71.110 396.170 ;
        RECT 71.950 395.720 73.870 396.170 ;
        RECT 74.710 395.720 76.630 396.170 ;
        RECT 77.470 395.720 79.390 396.170 ;
        RECT 80.230 395.720 82.150 396.170 ;
        RECT 82.990 395.720 84.910 396.170 ;
        RECT 85.750 395.720 87.670 396.170 ;
        RECT 88.510 395.720 90.430 396.170 ;
        RECT 91.270 395.720 93.190 396.170 ;
        RECT 94.030 395.720 95.950 396.170 ;
        RECT 96.790 395.720 98.710 396.170 ;
        RECT 99.550 395.720 101.470 396.170 ;
        RECT 102.310 395.720 104.230 396.170 ;
        RECT 105.070 395.720 106.990 396.170 ;
        RECT 107.830 395.720 109.750 396.170 ;
        RECT 110.590 395.720 112.510 396.170 ;
        RECT 113.350 395.720 115.270 396.170 ;
        RECT 116.110 395.720 118.030 396.170 ;
        RECT 118.870 395.720 120.790 396.170 ;
        RECT 121.630 395.720 123.550 396.170 ;
        RECT 124.390 395.720 126.310 396.170 ;
        RECT 127.150 395.720 129.070 396.170 ;
        RECT 129.910 395.720 131.830 396.170 ;
        RECT 132.670 395.720 134.590 396.170 ;
        RECT 135.430 395.720 137.350 396.170 ;
        RECT 138.190 395.720 140.110 396.170 ;
        RECT 140.950 395.720 142.870 396.170 ;
        RECT 143.710 395.720 145.630 396.170 ;
        RECT 146.470 395.720 148.390 396.170 ;
        RECT 149.230 395.720 151.150 396.170 ;
        RECT 151.990 395.720 153.910 396.170 ;
        RECT 154.750 395.720 156.670 396.170 ;
        RECT 157.510 395.720 159.430 396.170 ;
        RECT 160.270 395.720 162.190 396.170 ;
        RECT 163.030 395.720 164.950 396.170 ;
        RECT 165.790 395.720 167.710 396.170 ;
        RECT 168.550 395.720 170.470 396.170 ;
        RECT 171.310 395.720 173.230 396.170 ;
        RECT 174.070 395.720 175.990 396.170 ;
        RECT 176.830 395.720 178.750 396.170 ;
        RECT 179.590 395.720 181.510 396.170 ;
        RECT 182.350 395.720 184.270 396.170 ;
        RECT 185.110 395.720 187.030 396.170 ;
        RECT 187.870 395.720 189.790 396.170 ;
        RECT 190.630 395.720 192.550 396.170 ;
        RECT 193.390 395.720 195.310 396.170 ;
        RECT 196.150 395.720 198.070 396.170 ;
        RECT 198.910 395.720 200.830 396.170 ;
        RECT 201.670 395.720 203.590 396.170 ;
        RECT 204.430 395.720 206.350 396.170 ;
        RECT 207.190 395.720 209.110 396.170 ;
        RECT 209.950 395.720 211.870 396.170 ;
        RECT 212.710 395.720 214.630 396.170 ;
        RECT 215.470 395.720 217.390 396.170 ;
        RECT 218.230 395.720 220.150 396.170 ;
        RECT 220.990 395.720 222.910 396.170 ;
        RECT 223.750 395.720 225.670 396.170 ;
        RECT 226.510 395.720 228.430 396.170 ;
        RECT 229.270 395.720 231.190 396.170 ;
        RECT 232.030 395.720 233.950 396.170 ;
        RECT 234.790 395.720 236.710 396.170 ;
        RECT 237.550 395.720 239.470 396.170 ;
        RECT 240.310 395.720 242.230 396.170 ;
        RECT 243.070 395.720 244.990 396.170 ;
        RECT 245.830 395.720 247.750 396.170 ;
        RECT 248.590 395.720 250.510 396.170 ;
        RECT 251.350 395.720 253.270 396.170 ;
        RECT 254.110 395.720 256.030 396.170 ;
        RECT 256.870 395.720 258.790 396.170 ;
        RECT 259.630 395.720 261.550 396.170 ;
        RECT 262.390 395.720 264.310 396.170 ;
        RECT 265.150 395.720 267.070 396.170 ;
        RECT 267.910 395.720 269.830 396.170 ;
        RECT 270.670 395.720 272.590 396.170 ;
        RECT 273.430 395.720 275.350 396.170 ;
        RECT 276.190 395.720 278.110 396.170 ;
        RECT 278.950 395.720 280.870 396.170 ;
        RECT 281.710 395.720 283.630 396.170 ;
        RECT 284.470 395.720 286.390 396.170 ;
        RECT 287.230 395.720 289.150 396.170 ;
        RECT 289.990 395.720 291.910 396.170 ;
        RECT 292.750 395.720 294.670 396.170 ;
        RECT 295.510 395.720 297.430 396.170 ;
        RECT 298.270 395.720 300.190 396.170 ;
        RECT 301.030 395.720 302.950 396.170 ;
        RECT 303.790 395.720 305.710 396.170 ;
        RECT 306.550 395.720 308.470 396.170 ;
        RECT 309.310 395.720 311.230 396.170 ;
        RECT 312.070 395.720 313.990 396.170 ;
        RECT 314.830 395.720 316.750 396.170 ;
        RECT 317.590 395.720 319.510 396.170 ;
        RECT 320.350 395.720 322.270 396.170 ;
        RECT 323.110 395.720 325.030 396.170 ;
        RECT 325.870 395.720 327.790 396.170 ;
        RECT 328.630 395.720 330.550 396.170 ;
        RECT 331.390 395.720 333.310 396.170 ;
        RECT 334.150 395.720 336.070 396.170 ;
        RECT 336.910 395.720 338.830 396.170 ;
        RECT 339.670 395.720 341.590 396.170 ;
        RECT 342.430 395.720 344.350 396.170 ;
        RECT 345.190 395.720 347.110 396.170 ;
        RECT 347.950 395.720 349.870 396.170 ;
        RECT 350.710 395.720 352.630 396.170 ;
        RECT 353.470 395.720 355.390 396.170 ;
        RECT 356.230 395.720 358.150 396.170 ;
        RECT 358.990 395.720 360.910 396.170 ;
        RECT 361.750 395.720 363.670 396.170 ;
        RECT 364.510 395.720 366.430 396.170 ;
        RECT 367.270 395.720 369.190 396.170 ;
        RECT 370.030 395.720 371.950 396.170 ;
        RECT 372.790 395.720 374.710 396.170 ;
        RECT 375.550 395.720 377.470 396.170 ;
        RECT 378.310 395.720 380.230 396.170 ;
        RECT 381.070 395.720 382.990 396.170 ;
        RECT 383.830 395.720 385.750 396.170 ;
        RECT 386.590 395.720 388.510 396.170 ;
        RECT 389.350 395.720 395.510 396.170 ;
        RECT 4.690 4.280 395.510 395.720 ;
        RECT 4.690 1.515 14.530 4.280 ;
        RECT 15.370 1.515 20.050 4.280 ;
        RECT 20.890 1.515 25.570 4.280 ;
        RECT 26.410 1.515 31.090 4.280 ;
        RECT 31.930 1.515 36.610 4.280 ;
        RECT 37.450 1.515 42.130 4.280 ;
        RECT 42.970 1.515 47.650 4.280 ;
        RECT 48.490 1.515 53.170 4.280 ;
        RECT 54.010 1.515 58.690 4.280 ;
        RECT 59.530 1.515 64.210 4.280 ;
        RECT 65.050 1.515 69.730 4.280 ;
        RECT 70.570 1.515 75.250 4.280 ;
        RECT 76.090 1.515 80.770 4.280 ;
        RECT 81.610 1.515 86.290 4.280 ;
        RECT 87.130 1.515 91.810 4.280 ;
        RECT 92.650 1.515 97.330 4.280 ;
        RECT 98.170 1.515 102.850 4.280 ;
        RECT 103.690 1.515 108.370 4.280 ;
        RECT 109.210 1.515 113.890 4.280 ;
        RECT 114.730 1.515 119.410 4.280 ;
        RECT 120.250 1.515 124.930 4.280 ;
        RECT 125.770 1.515 130.450 4.280 ;
        RECT 131.290 1.515 135.970 4.280 ;
        RECT 136.810 1.515 141.490 4.280 ;
        RECT 142.330 1.515 147.010 4.280 ;
        RECT 147.850 1.515 152.530 4.280 ;
        RECT 153.370 1.515 158.050 4.280 ;
        RECT 158.890 1.515 163.570 4.280 ;
        RECT 164.410 1.515 169.090 4.280 ;
        RECT 169.930 1.515 174.610 4.280 ;
        RECT 175.450 1.515 180.130 4.280 ;
        RECT 180.970 1.515 185.650 4.280 ;
        RECT 186.490 1.515 191.170 4.280 ;
        RECT 192.010 1.515 196.690 4.280 ;
        RECT 197.530 1.515 202.210 4.280 ;
        RECT 203.050 1.515 207.730 4.280 ;
        RECT 208.570 1.515 213.250 4.280 ;
        RECT 214.090 1.515 218.770 4.280 ;
        RECT 219.610 1.515 224.290 4.280 ;
        RECT 225.130 1.515 229.810 4.280 ;
        RECT 230.650 1.515 235.330 4.280 ;
        RECT 236.170 1.515 240.850 4.280 ;
        RECT 241.690 1.515 246.370 4.280 ;
        RECT 247.210 1.515 251.890 4.280 ;
        RECT 252.730 1.515 257.410 4.280 ;
        RECT 258.250 1.515 262.930 4.280 ;
        RECT 263.770 1.515 268.450 4.280 ;
        RECT 269.290 1.515 273.970 4.280 ;
        RECT 274.810 1.515 279.490 4.280 ;
        RECT 280.330 1.515 285.010 4.280 ;
        RECT 285.850 1.515 290.530 4.280 ;
        RECT 291.370 1.515 296.050 4.280 ;
        RECT 296.890 1.515 301.570 4.280 ;
        RECT 302.410 1.515 307.090 4.280 ;
        RECT 307.930 1.515 312.610 4.280 ;
        RECT 313.450 1.515 318.130 4.280 ;
        RECT 318.970 1.515 323.650 4.280 ;
        RECT 324.490 1.515 329.170 4.280 ;
        RECT 330.010 1.515 334.690 4.280 ;
        RECT 335.530 1.515 340.210 4.280 ;
        RECT 341.050 1.515 345.730 4.280 ;
        RECT 346.570 1.515 351.250 4.280 ;
        RECT 352.090 1.515 356.770 4.280 ;
        RECT 357.610 1.515 362.290 4.280 ;
        RECT 363.130 1.515 367.810 4.280 ;
        RECT 368.650 1.515 373.330 4.280 ;
        RECT 374.170 1.515 378.850 4.280 ;
        RECT 379.690 1.515 384.370 4.280 ;
        RECT 385.210 1.515 395.510 4.280 ;
      LAYER met3 ;
        RECT 4.400 396.760 396.000 397.610 ;
        RECT 3.990 394.080 396.000 396.760 ;
        RECT 4.400 392.680 396.000 394.080 ;
        RECT 3.990 390.000 396.000 392.680 ;
        RECT 4.400 388.600 396.000 390.000 ;
        RECT 3.990 385.920 396.000 388.600 ;
        RECT 4.400 384.520 396.000 385.920 ;
        RECT 3.990 381.840 396.000 384.520 ;
        RECT 4.400 380.440 396.000 381.840 ;
        RECT 3.990 377.760 396.000 380.440 ;
        RECT 4.400 376.360 396.000 377.760 ;
        RECT 3.990 373.680 396.000 376.360 ;
        RECT 4.400 372.280 396.000 373.680 ;
        RECT 3.990 369.600 396.000 372.280 ;
        RECT 4.400 368.200 396.000 369.600 ;
        RECT 3.990 365.520 396.000 368.200 ;
        RECT 4.400 364.120 396.000 365.520 ;
        RECT 3.990 361.440 396.000 364.120 ;
        RECT 4.400 360.040 396.000 361.440 ;
        RECT 3.990 357.360 396.000 360.040 ;
        RECT 4.400 355.960 396.000 357.360 ;
        RECT 3.990 353.280 396.000 355.960 ;
        RECT 4.400 351.880 396.000 353.280 ;
        RECT 3.990 349.200 396.000 351.880 ;
        RECT 4.400 347.800 396.000 349.200 ;
        RECT 3.990 345.120 396.000 347.800 ;
        RECT 4.400 343.720 395.600 345.120 ;
        RECT 3.990 342.400 396.000 343.720 ;
        RECT 3.990 341.040 395.600 342.400 ;
        RECT 4.400 341.000 395.600 341.040 ;
        RECT 4.400 339.680 396.000 341.000 ;
        RECT 4.400 339.640 395.600 339.680 ;
        RECT 3.990 338.280 395.600 339.640 ;
        RECT 3.990 336.960 396.000 338.280 ;
        RECT 4.400 335.560 395.600 336.960 ;
        RECT 3.990 334.240 396.000 335.560 ;
        RECT 3.990 332.880 395.600 334.240 ;
        RECT 4.400 332.840 395.600 332.880 ;
        RECT 4.400 331.520 396.000 332.840 ;
        RECT 4.400 331.480 395.600 331.520 ;
        RECT 3.990 330.120 395.600 331.480 ;
        RECT 3.990 328.800 396.000 330.120 ;
        RECT 4.400 327.400 395.600 328.800 ;
        RECT 3.990 326.080 396.000 327.400 ;
        RECT 3.990 324.720 395.600 326.080 ;
        RECT 4.400 324.680 395.600 324.720 ;
        RECT 4.400 323.360 396.000 324.680 ;
        RECT 4.400 323.320 395.600 323.360 ;
        RECT 3.990 321.960 395.600 323.320 ;
        RECT 3.990 320.640 396.000 321.960 ;
        RECT 4.400 319.240 395.600 320.640 ;
        RECT 3.990 317.920 396.000 319.240 ;
        RECT 3.990 316.560 395.600 317.920 ;
        RECT 4.400 316.520 395.600 316.560 ;
        RECT 4.400 315.200 396.000 316.520 ;
        RECT 4.400 315.160 395.600 315.200 ;
        RECT 3.990 313.800 395.600 315.160 ;
        RECT 3.990 312.480 396.000 313.800 ;
        RECT 4.400 311.080 395.600 312.480 ;
        RECT 3.990 309.760 396.000 311.080 ;
        RECT 3.990 308.400 395.600 309.760 ;
        RECT 4.400 308.360 395.600 308.400 ;
        RECT 4.400 307.040 396.000 308.360 ;
        RECT 4.400 307.000 395.600 307.040 ;
        RECT 3.990 305.640 395.600 307.000 ;
        RECT 3.990 304.320 396.000 305.640 ;
        RECT 4.400 302.920 395.600 304.320 ;
        RECT 3.990 301.600 396.000 302.920 ;
        RECT 3.990 300.240 395.600 301.600 ;
        RECT 4.400 300.200 395.600 300.240 ;
        RECT 4.400 298.880 396.000 300.200 ;
        RECT 4.400 298.840 395.600 298.880 ;
        RECT 3.990 297.480 395.600 298.840 ;
        RECT 3.990 296.160 396.000 297.480 ;
        RECT 4.400 294.760 395.600 296.160 ;
        RECT 3.990 293.440 396.000 294.760 ;
        RECT 3.990 292.080 395.600 293.440 ;
        RECT 4.400 292.040 395.600 292.080 ;
        RECT 4.400 290.720 396.000 292.040 ;
        RECT 4.400 290.680 395.600 290.720 ;
        RECT 3.990 289.320 395.600 290.680 ;
        RECT 3.990 288.000 396.000 289.320 ;
        RECT 4.400 286.600 395.600 288.000 ;
        RECT 3.990 285.280 396.000 286.600 ;
        RECT 3.990 283.920 395.600 285.280 ;
        RECT 4.400 283.880 395.600 283.920 ;
        RECT 4.400 282.560 396.000 283.880 ;
        RECT 4.400 282.520 395.600 282.560 ;
        RECT 3.990 281.160 395.600 282.520 ;
        RECT 3.990 279.840 396.000 281.160 ;
        RECT 4.400 278.440 395.600 279.840 ;
        RECT 3.990 277.120 396.000 278.440 ;
        RECT 3.990 275.760 395.600 277.120 ;
        RECT 4.400 275.720 395.600 275.760 ;
        RECT 4.400 274.400 396.000 275.720 ;
        RECT 4.400 274.360 395.600 274.400 ;
        RECT 3.990 273.000 395.600 274.360 ;
        RECT 3.990 271.680 396.000 273.000 ;
        RECT 4.400 270.280 395.600 271.680 ;
        RECT 3.990 268.960 396.000 270.280 ;
        RECT 3.990 267.600 395.600 268.960 ;
        RECT 4.400 267.560 395.600 267.600 ;
        RECT 4.400 266.240 396.000 267.560 ;
        RECT 4.400 266.200 395.600 266.240 ;
        RECT 3.990 264.840 395.600 266.200 ;
        RECT 3.990 263.520 396.000 264.840 ;
        RECT 4.400 262.120 395.600 263.520 ;
        RECT 3.990 260.800 396.000 262.120 ;
        RECT 3.990 259.440 395.600 260.800 ;
        RECT 4.400 259.400 395.600 259.440 ;
        RECT 4.400 258.080 396.000 259.400 ;
        RECT 4.400 258.040 395.600 258.080 ;
        RECT 3.990 256.680 395.600 258.040 ;
        RECT 3.990 255.360 396.000 256.680 ;
        RECT 4.400 253.960 395.600 255.360 ;
        RECT 3.990 252.640 396.000 253.960 ;
        RECT 3.990 251.280 395.600 252.640 ;
        RECT 4.400 251.240 395.600 251.280 ;
        RECT 4.400 249.920 396.000 251.240 ;
        RECT 4.400 249.880 395.600 249.920 ;
        RECT 3.990 248.520 395.600 249.880 ;
        RECT 3.990 247.200 396.000 248.520 ;
        RECT 4.400 245.800 395.600 247.200 ;
        RECT 3.990 244.480 396.000 245.800 ;
        RECT 3.990 243.120 395.600 244.480 ;
        RECT 4.400 243.080 395.600 243.120 ;
        RECT 4.400 241.760 396.000 243.080 ;
        RECT 4.400 241.720 395.600 241.760 ;
        RECT 3.990 240.360 395.600 241.720 ;
        RECT 3.990 239.040 396.000 240.360 ;
        RECT 4.400 237.640 395.600 239.040 ;
        RECT 3.990 236.320 396.000 237.640 ;
        RECT 3.990 234.960 395.600 236.320 ;
        RECT 4.400 234.920 395.600 234.960 ;
        RECT 4.400 233.600 396.000 234.920 ;
        RECT 4.400 233.560 395.600 233.600 ;
        RECT 3.990 232.200 395.600 233.560 ;
        RECT 3.990 230.880 396.000 232.200 ;
        RECT 4.400 229.480 395.600 230.880 ;
        RECT 3.990 228.160 396.000 229.480 ;
        RECT 3.990 226.800 395.600 228.160 ;
        RECT 4.400 226.760 395.600 226.800 ;
        RECT 4.400 225.440 396.000 226.760 ;
        RECT 4.400 225.400 395.600 225.440 ;
        RECT 3.990 224.040 395.600 225.400 ;
        RECT 3.990 222.720 396.000 224.040 ;
        RECT 4.400 221.320 395.600 222.720 ;
        RECT 3.990 220.000 396.000 221.320 ;
        RECT 3.990 218.640 395.600 220.000 ;
        RECT 4.400 218.600 395.600 218.640 ;
        RECT 4.400 217.280 396.000 218.600 ;
        RECT 4.400 217.240 395.600 217.280 ;
        RECT 3.990 215.880 395.600 217.240 ;
        RECT 3.990 214.560 396.000 215.880 ;
        RECT 4.400 213.160 395.600 214.560 ;
        RECT 3.990 211.840 396.000 213.160 ;
        RECT 3.990 210.480 395.600 211.840 ;
        RECT 4.400 210.440 395.600 210.480 ;
        RECT 4.400 209.120 396.000 210.440 ;
        RECT 4.400 209.080 395.600 209.120 ;
        RECT 3.990 207.720 395.600 209.080 ;
        RECT 3.990 206.400 396.000 207.720 ;
        RECT 4.400 205.000 395.600 206.400 ;
        RECT 3.990 203.680 396.000 205.000 ;
        RECT 3.990 202.320 395.600 203.680 ;
        RECT 4.400 202.280 395.600 202.320 ;
        RECT 4.400 200.960 396.000 202.280 ;
        RECT 4.400 200.920 395.600 200.960 ;
        RECT 3.990 199.560 395.600 200.920 ;
        RECT 3.990 198.240 396.000 199.560 ;
        RECT 4.400 196.840 395.600 198.240 ;
        RECT 3.990 195.520 396.000 196.840 ;
        RECT 3.990 194.160 395.600 195.520 ;
        RECT 4.400 194.120 395.600 194.160 ;
        RECT 4.400 192.800 396.000 194.120 ;
        RECT 4.400 192.760 395.600 192.800 ;
        RECT 3.990 191.400 395.600 192.760 ;
        RECT 3.990 190.080 396.000 191.400 ;
        RECT 4.400 188.680 395.600 190.080 ;
        RECT 3.990 187.360 396.000 188.680 ;
        RECT 3.990 186.000 395.600 187.360 ;
        RECT 4.400 185.960 395.600 186.000 ;
        RECT 4.400 184.640 396.000 185.960 ;
        RECT 4.400 184.600 395.600 184.640 ;
        RECT 3.990 183.240 395.600 184.600 ;
        RECT 3.990 181.920 396.000 183.240 ;
        RECT 4.400 180.520 395.600 181.920 ;
        RECT 3.990 179.200 396.000 180.520 ;
        RECT 3.990 177.840 395.600 179.200 ;
        RECT 4.400 177.800 395.600 177.840 ;
        RECT 4.400 176.480 396.000 177.800 ;
        RECT 4.400 176.440 395.600 176.480 ;
        RECT 3.990 175.080 395.600 176.440 ;
        RECT 3.990 173.760 396.000 175.080 ;
        RECT 4.400 172.360 395.600 173.760 ;
        RECT 3.990 171.040 396.000 172.360 ;
        RECT 3.990 169.680 395.600 171.040 ;
        RECT 4.400 169.640 395.600 169.680 ;
        RECT 4.400 168.320 396.000 169.640 ;
        RECT 4.400 168.280 395.600 168.320 ;
        RECT 3.990 166.920 395.600 168.280 ;
        RECT 3.990 165.600 396.000 166.920 ;
        RECT 4.400 164.200 395.600 165.600 ;
        RECT 3.990 162.880 396.000 164.200 ;
        RECT 3.990 161.520 395.600 162.880 ;
        RECT 4.400 161.480 395.600 161.520 ;
        RECT 4.400 160.160 396.000 161.480 ;
        RECT 4.400 160.120 395.600 160.160 ;
        RECT 3.990 158.760 395.600 160.120 ;
        RECT 3.990 157.440 396.000 158.760 ;
        RECT 4.400 156.040 395.600 157.440 ;
        RECT 3.990 154.720 396.000 156.040 ;
        RECT 3.990 153.360 395.600 154.720 ;
        RECT 4.400 153.320 395.600 153.360 ;
        RECT 4.400 152.000 396.000 153.320 ;
        RECT 4.400 151.960 395.600 152.000 ;
        RECT 3.990 150.600 395.600 151.960 ;
        RECT 3.990 149.280 396.000 150.600 ;
        RECT 4.400 147.880 395.600 149.280 ;
        RECT 3.990 146.560 396.000 147.880 ;
        RECT 3.990 145.200 395.600 146.560 ;
        RECT 4.400 145.160 395.600 145.200 ;
        RECT 4.400 143.840 396.000 145.160 ;
        RECT 4.400 143.800 395.600 143.840 ;
        RECT 3.990 142.440 395.600 143.800 ;
        RECT 3.990 141.120 396.000 142.440 ;
        RECT 4.400 139.720 395.600 141.120 ;
        RECT 3.990 138.400 396.000 139.720 ;
        RECT 3.990 137.040 395.600 138.400 ;
        RECT 4.400 137.000 395.600 137.040 ;
        RECT 4.400 135.680 396.000 137.000 ;
        RECT 4.400 135.640 395.600 135.680 ;
        RECT 3.990 134.280 395.600 135.640 ;
        RECT 3.990 132.960 396.000 134.280 ;
        RECT 4.400 131.560 395.600 132.960 ;
        RECT 3.990 130.240 396.000 131.560 ;
        RECT 3.990 128.880 395.600 130.240 ;
        RECT 4.400 128.840 395.600 128.880 ;
        RECT 4.400 127.520 396.000 128.840 ;
        RECT 4.400 127.480 395.600 127.520 ;
        RECT 3.990 126.120 395.600 127.480 ;
        RECT 3.990 124.800 396.000 126.120 ;
        RECT 4.400 123.400 395.600 124.800 ;
        RECT 3.990 122.080 396.000 123.400 ;
        RECT 3.990 120.720 395.600 122.080 ;
        RECT 4.400 120.680 395.600 120.720 ;
        RECT 4.400 119.360 396.000 120.680 ;
        RECT 4.400 119.320 395.600 119.360 ;
        RECT 3.990 117.960 395.600 119.320 ;
        RECT 3.990 116.640 396.000 117.960 ;
        RECT 4.400 115.240 395.600 116.640 ;
        RECT 3.990 113.920 396.000 115.240 ;
        RECT 3.990 112.560 395.600 113.920 ;
        RECT 4.400 112.520 395.600 112.560 ;
        RECT 4.400 111.200 396.000 112.520 ;
        RECT 4.400 111.160 395.600 111.200 ;
        RECT 3.990 109.800 395.600 111.160 ;
        RECT 3.990 108.480 396.000 109.800 ;
        RECT 4.400 107.080 395.600 108.480 ;
        RECT 3.990 105.760 396.000 107.080 ;
        RECT 3.990 104.400 395.600 105.760 ;
        RECT 4.400 104.360 395.600 104.400 ;
        RECT 4.400 103.040 396.000 104.360 ;
        RECT 4.400 103.000 395.600 103.040 ;
        RECT 3.990 101.640 395.600 103.000 ;
        RECT 3.990 100.320 396.000 101.640 ;
        RECT 4.400 98.920 395.600 100.320 ;
        RECT 3.990 97.600 396.000 98.920 ;
        RECT 3.990 96.240 395.600 97.600 ;
        RECT 4.400 96.200 395.600 96.240 ;
        RECT 4.400 94.880 396.000 96.200 ;
        RECT 4.400 94.840 395.600 94.880 ;
        RECT 3.990 93.480 395.600 94.840 ;
        RECT 3.990 92.160 396.000 93.480 ;
        RECT 4.400 90.760 395.600 92.160 ;
        RECT 3.990 89.440 396.000 90.760 ;
        RECT 3.990 88.080 395.600 89.440 ;
        RECT 4.400 88.040 395.600 88.080 ;
        RECT 4.400 86.720 396.000 88.040 ;
        RECT 4.400 86.680 395.600 86.720 ;
        RECT 3.990 85.320 395.600 86.680 ;
        RECT 3.990 84.000 396.000 85.320 ;
        RECT 4.400 82.600 395.600 84.000 ;
        RECT 3.990 81.280 396.000 82.600 ;
        RECT 3.990 79.920 395.600 81.280 ;
        RECT 4.400 79.880 395.600 79.920 ;
        RECT 4.400 78.560 396.000 79.880 ;
        RECT 4.400 78.520 395.600 78.560 ;
        RECT 3.990 77.160 395.600 78.520 ;
        RECT 3.990 75.840 396.000 77.160 ;
        RECT 4.400 74.440 395.600 75.840 ;
        RECT 3.990 73.120 396.000 74.440 ;
        RECT 3.990 71.760 395.600 73.120 ;
        RECT 4.400 71.720 395.600 71.760 ;
        RECT 4.400 70.400 396.000 71.720 ;
        RECT 4.400 70.360 395.600 70.400 ;
        RECT 3.990 69.000 395.600 70.360 ;
        RECT 3.990 67.680 396.000 69.000 ;
        RECT 4.400 66.280 395.600 67.680 ;
        RECT 3.990 64.960 396.000 66.280 ;
        RECT 3.990 63.600 395.600 64.960 ;
        RECT 4.400 63.560 395.600 63.600 ;
        RECT 4.400 62.240 396.000 63.560 ;
        RECT 4.400 62.200 395.600 62.240 ;
        RECT 3.990 60.840 395.600 62.200 ;
        RECT 3.990 59.520 396.000 60.840 ;
        RECT 4.400 58.120 395.600 59.520 ;
        RECT 3.990 56.800 396.000 58.120 ;
        RECT 3.990 55.440 395.600 56.800 ;
        RECT 4.400 55.400 395.600 55.440 ;
        RECT 4.400 54.080 396.000 55.400 ;
        RECT 4.400 54.040 395.600 54.080 ;
        RECT 3.990 52.680 395.600 54.040 ;
        RECT 3.990 51.360 396.000 52.680 ;
        RECT 4.400 49.960 396.000 51.360 ;
        RECT 3.990 47.280 396.000 49.960 ;
        RECT 4.400 45.880 396.000 47.280 ;
        RECT 3.990 43.200 396.000 45.880 ;
        RECT 4.400 41.800 396.000 43.200 ;
        RECT 3.990 39.120 396.000 41.800 ;
        RECT 4.400 37.720 396.000 39.120 ;
        RECT 3.990 35.040 396.000 37.720 ;
        RECT 4.400 33.640 396.000 35.040 ;
        RECT 3.990 30.960 396.000 33.640 ;
        RECT 4.400 29.560 396.000 30.960 ;
        RECT 3.990 26.880 396.000 29.560 ;
        RECT 4.400 25.480 396.000 26.880 ;
        RECT 3.990 22.800 396.000 25.480 ;
        RECT 4.400 21.400 396.000 22.800 ;
        RECT 3.990 18.720 396.000 21.400 ;
        RECT 4.400 17.320 396.000 18.720 ;
        RECT 3.990 14.640 396.000 17.320 ;
        RECT 4.400 13.240 396.000 14.640 ;
        RECT 3.990 10.560 396.000 13.240 ;
        RECT 4.400 9.160 396.000 10.560 ;
        RECT 3.990 6.480 396.000 9.160 ;
        RECT 4.400 5.080 396.000 6.480 ;
        RECT 3.990 2.400 396.000 5.080 ;
        RECT 4.400 1.535 396.000 2.400 ;
      LAYER met4 ;
        RECT 25.135 96.055 97.440 379.945 ;
        RECT 99.840 96.055 174.240 379.945 ;
        RECT 176.640 96.055 230.625 379.945 ;
  END
END datapath
END LIBRARY

