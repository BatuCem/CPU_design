VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO registerFile
  CLASS BLOCK ;
  FOREIGN registerFile ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END clk
  PIN readAddr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END readAddr1[0]
  PIN readAddr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END readAddr1[1]
  PIN readAddr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END readAddr1[2]
  PIN readAddr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END readAddr1[3]
  PIN readAddr1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END readAddr1[4]
  PIN readAddr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END readAddr2[0]
  PIN readAddr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END readAddr2[1]
  PIN readAddr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END readAddr2[2]
  PIN readAddr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END readAddr2[3]
  PIN readAddr2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END readAddr2[4]
  PIN readData1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END readData1[0]
  PIN readData1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END readData1[10]
  PIN readData1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END readData1[11]
  PIN readData1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END readData1[12]
  PIN readData1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END readData1[13]
  PIN readData1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END readData1[14]
  PIN readData1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END readData1[15]
  PIN readData1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END readData1[16]
  PIN readData1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END readData1[17]
  PIN readData1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END readData1[18]
  PIN readData1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END readData1[19]
  PIN readData1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END readData1[1]
  PIN readData1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END readData1[20]
  PIN readData1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END readData1[21]
  PIN readData1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END readData1[22]
  PIN readData1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END readData1[23]
  PIN readData1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END readData1[24]
  PIN readData1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END readData1[25]
  PIN readData1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END readData1[26]
  PIN readData1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END readData1[27]
  PIN readData1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END readData1[28]
  PIN readData1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END readData1[29]
  PIN readData1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END readData1[2]
  PIN readData1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END readData1[30]
  PIN readData1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END readData1[31]
  PIN readData1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END readData1[3]
  PIN readData1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END readData1[4]
  PIN readData1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END readData1[5]
  PIN readData1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END readData1[6]
  PIN readData1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END readData1[7]
  PIN readData1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END readData1[8]
  PIN readData1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END readData1[9]
  PIN readData2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END readData2[0]
  PIN readData2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END readData2[10]
  PIN readData2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END readData2[11]
  PIN readData2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END readData2[12]
  PIN readData2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END readData2[13]
  PIN readData2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END readData2[14]
  PIN readData2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END readData2[15]
  PIN readData2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END readData2[16]
  PIN readData2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END readData2[17]
  PIN readData2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END readData2[18]
  PIN readData2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END readData2[19]
  PIN readData2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END readData2[1]
  PIN readData2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END readData2[20]
  PIN readData2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END readData2[21]
  PIN readData2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END readData2[22]
  PIN readData2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END readData2[23]
  PIN readData2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END readData2[24]
  PIN readData2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END readData2[25]
  PIN readData2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END readData2[26]
  PIN readData2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END readData2[27]
  PIN readData2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END readData2[28]
  PIN readData2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END readData2[29]
  PIN readData2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END readData2[2]
  PIN readData2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END readData2[30]
  PIN readData2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END readData2[31]
  PIN readData2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END readData2[3]
  PIN readData2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END readData2[4]
  PIN readData2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END readData2[5]
  PIN readData2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END readData2[6]
  PIN readData2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END readData2[7]
  PIN readData2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END readData2[8]
  PIN readData2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END readData2[9]
  PIN writeAddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END writeAddr[0]
  PIN writeAddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END writeAddr[1]
  PIN writeAddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END writeAddr[2]
  PIN writeAddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END writeAddr[3]
  PIN writeAddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END writeAddr[4]
  PIN writeData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END writeData[0]
  PIN writeData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END writeData[10]
  PIN writeData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END writeData[11]
  PIN writeData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END writeData[12]
  PIN writeData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END writeData[13]
  PIN writeData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END writeData[14]
  PIN writeData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END writeData[15]
  PIN writeData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END writeData[16]
  PIN writeData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END writeData[17]
  PIN writeData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END writeData[18]
  PIN writeData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END writeData[19]
  PIN writeData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END writeData[1]
  PIN writeData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END writeData[20]
  PIN writeData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END writeData[21]
  PIN writeData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END writeData[22]
  PIN writeData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END writeData[23]
  PIN writeData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END writeData[24]
  PIN writeData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END writeData[25]
  PIN writeData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END writeData[26]
  PIN writeData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END writeData[27]
  PIN writeData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END writeData[28]
  PIN writeData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END writeData[29]
  PIN writeData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END writeData[2]
  PIN writeData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END writeData[30]
  PIN writeData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END writeData[31]
  PIN writeData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END writeData[3]
  PIN writeData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END writeData[4]
  PIN writeData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END writeData[5]
  PIN writeData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END writeData[6]
  PIN writeData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END writeData[7]
  PIN writeData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END writeData[8]
  PIN writeData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END writeData[9]
  PIN writeEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END writeEn
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 587.605 ;
      LAYER met1 ;
        RECT 4.670 10.640 594.620 587.760 ;
      LAYER met2 ;
        RECT 4.690 10.695 592.840 587.705 ;
      LAYER met3 ;
        RECT 3.990 528.720 574.475 587.685 ;
        RECT 4.400 527.320 574.475 528.720 ;
        RECT 3.990 524.640 574.475 527.320 ;
        RECT 4.400 523.240 574.475 524.640 ;
        RECT 3.990 520.560 574.475 523.240 ;
        RECT 4.400 519.160 574.475 520.560 ;
        RECT 3.990 516.480 574.475 519.160 ;
        RECT 4.400 515.080 574.475 516.480 ;
        RECT 3.990 512.400 574.475 515.080 ;
        RECT 4.400 511.000 574.475 512.400 ;
        RECT 3.990 508.320 574.475 511.000 ;
        RECT 4.400 506.920 574.475 508.320 ;
        RECT 3.990 504.240 574.475 506.920 ;
        RECT 4.400 502.840 574.475 504.240 ;
        RECT 3.990 500.160 574.475 502.840 ;
        RECT 4.400 498.760 574.475 500.160 ;
        RECT 3.990 496.080 574.475 498.760 ;
        RECT 4.400 494.680 574.475 496.080 ;
        RECT 3.990 492.000 574.475 494.680 ;
        RECT 4.400 490.600 574.475 492.000 ;
        RECT 3.990 487.920 574.475 490.600 ;
        RECT 4.400 486.520 574.475 487.920 ;
        RECT 3.990 483.840 574.475 486.520 ;
        RECT 4.400 482.440 574.475 483.840 ;
        RECT 3.990 479.760 574.475 482.440 ;
        RECT 4.400 478.360 574.475 479.760 ;
        RECT 3.990 475.680 574.475 478.360 ;
        RECT 4.400 474.280 574.475 475.680 ;
        RECT 3.990 471.600 574.475 474.280 ;
        RECT 4.400 470.200 574.475 471.600 ;
        RECT 3.990 467.520 574.475 470.200 ;
        RECT 4.400 466.120 574.475 467.520 ;
        RECT 3.990 463.440 574.475 466.120 ;
        RECT 4.400 462.040 574.475 463.440 ;
        RECT 3.990 459.360 574.475 462.040 ;
        RECT 4.400 457.960 574.475 459.360 ;
        RECT 3.990 455.280 574.475 457.960 ;
        RECT 4.400 453.880 574.475 455.280 ;
        RECT 3.990 451.200 574.475 453.880 ;
        RECT 4.400 449.800 574.475 451.200 ;
        RECT 3.990 447.120 574.475 449.800 ;
        RECT 4.400 445.720 574.475 447.120 ;
        RECT 3.990 443.040 574.475 445.720 ;
        RECT 4.400 441.640 574.475 443.040 ;
        RECT 3.990 438.960 574.475 441.640 ;
        RECT 4.400 437.560 574.475 438.960 ;
        RECT 3.990 434.880 574.475 437.560 ;
        RECT 4.400 433.480 574.475 434.880 ;
        RECT 3.990 430.800 574.475 433.480 ;
        RECT 4.400 429.400 574.475 430.800 ;
        RECT 3.990 426.720 574.475 429.400 ;
        RECT 4.400 425.320 574.475 426.720 ;
        RECT 3.990 422.640 574.475 425.320 ;
        RECT 4.400 421.240 574.475 422.640 ;
        RECT 3.990 418.560 574.475 421.240 ;
        RECT 4.400 417.160 574.475 418.560 ;
        RECT 3.990 414.480 574.475 417.160 ;
        RECT 4.400 413.080 574.475 414.480 ;
        RECT 3.990 410.400 574.475 413.080 ;
        RECT 4.400 409.000 574.475 410.400 ;
        RECT 3.990 406.320 574.475 409.000 ;
        RECT 4.400 404.920 574.475 406.320 ;
        RECT 3.990 402.240 574.475 404.920 ;
        RECT 4.400 400.840 574.475 402.240 ;
        RECT 3.990 398.160 574.475 400.840 ;
        RECT 4.400 396.760 574.475 398.160 ;
        RECT 3.990 394.080 574.475 396.760 ;
        RECT 4.400 392.680 574.475 394.080 ;
        RECT 3.990 390.000 574.475 392.680 ;
        RECT 4.400 388.600 574.475 390.000 ;
        RECT 3.990 385.920 574.475 388.600 ;
        RECT 4.400 384.520 574.475 385.920 ;
        RECT 3.990 381.840 574.475 384.520 ;
        RECT 4.400 380.440 574.475 381.840 ;
        RECT 3.990 377.760 574.475 380.440 ;
        RECT 4.400 376.360 574.475 377.760 ;
        RECT 3.990 373.680 574.475 376.360 ;
        RECT 4.400 372.280 574.475 373.680 ;
        RECT 3.990 369.600 574.475 372.280 ;
        RECT 4.400 368.200 574.475 369.600 ;
        RECT 3.990 365.520 574.475 368.200 ;
        RECT 4.400 364.120 574.475 365.520 ;
        RECT 3.990 361.440 574.475 364.120 ;
        RECT 4.400 360.040 574.475 361.440 ;
        RECT 3.990 357.360 574.475 360.040 ;
        RECT 4.400 355.960 574.475 357.360 ;
        RECT 3.990 353.280 574.475 355.960 ;
        RECT 4.400 351.880 574.475 353.280 ;
        RECT 3.990 349.200 574.475 351.880 ;
        RECT 4.400 347.800 574.475 349.200 ;
        RECT 3.990 345.120 574.475 347.800 ;
        RECT 4.400 343.720 574.475 345.120 ;
        RECT 3.990 341.040 574.475 343.720 ;
        RECT 4.400 339.640 574.475 341.040 ;
        RECT 3.990 336.960 574.475 339.640 ;
        RECT 4.400 335.560 574.475 336.960 ;
        RECT 3.990 332.880 574.475 335.560 ;
        RECT 4.400 331.480 574.475 332.880 ;
        RECT 3.990 328.800 574.475 331.480 ;
        RECT 4.400 327.400 574.475 328.800 ;
        RECT 3.990 324.720 574.475 327.400 ;
        RECT 4.400 323.320 574.475 324.720 ;
        RECT 3.990 320.640 574.475 323.320 ;
        RECT 4.400 319.240 574.475 320.640 ;
        RECT 3.990 316.560 574.475 319.240 ;
        RECT 4.400 315.160 574.475 316.560 ;
        RECT 3.990 312.480 574.475 315.160 ;
        RECT 4.400 311.080 574.475 312.480 ;
        RECT 3.990 308.400 574.475 311.080 ;
        RECT 4.400 307.000 574.475 308.400 ;
        RECT 3.990 304.320 574.475 307.000 ;
        RECT 4.400 302.920 574.475 304.320 ;
        RECT 3.990 300.240 574.475 302.920 ;
        RECT 4.400 298.840 574.475 300.240 ;
        RECT 3.990 296.160 574.475 298.840 ;
        RECT 4.400 294.760 574.475 296.160 ;
        RECT 3.990 292.080 574.475 294.760 ;
        RECT 4.400 290.680 574.475 292.080 ;
        RECT 3.990 288.000 574.475 290.680 ;
        RECT 4.400 286.600 574.475 288.000 ;
        RECT 3.990 283.920 574.475 286.600 ;
        RECT 4.400 282.520 574.475 283.920 ;
        RECT 3.990 279.840 574.475 282.520 ;
        RECT 4.400 278.440 574.475 279.840 ;
        RECT 3.990 275.760 574.475 278.440 ;
        RECT 4.400 274.360 574.475 275.760 ;
        RECT 3.990 271.680 574.475 274.360 ;
        RECT 4.400 270.280 574.475 271.680 ;
        RECT 3.990 267.600 574.475 270.280 ;
        RECT 4.400 266.200 574.475 267.600 ;
        RECT 3.990 263.520 574.475 266.200 ;
        RECT 4.400 262.120 574.475 263.520 ;
        RECT 3.990 259.440 574.475 262.120 ;
        RECT 4.400 258.040 574.475 259.440 ;
        RECT 3.990 255.360 574.475 258.040 ;
        RECT 4.400 253.960 574.475 255.360 ;
        RECT 3.990 251.280 574.475 253.960 ;
        RECT 4.400 249.880 574.475 251.280 ;
        RECT 3.990 247.200 574.475 249.880 ;
        RECT 4.400 245.800 574.475 247.200 ;
        RECT 3.990 243.120 574.475 245.800 ;
        RECT 4.400 241.720 574.475 243.120 ;
        RECT 3.990 239.040 574.475 241.720 ;
        RECT 4.400 237.640 574.475 239.040 ;
        RECT 3.990 234.960 574.475 237.640 ;
        RECT 4.400 233.560 574.475 234.960 ;
        RECT 3.990 230.880 574.475 233.560 ;
        RECT 4.400 229.480 574.475 230.880 ;
        RECT 3.990 226.800 574.475 229.480 ;
        RECT 4.400 225.400 574.475 226.800 ;
        RECT 3.990 222.720 574.475 225.400 ;
        RECT 4.400 221.320 574.475 222.720 ;
        RECT 3.990 218.640 574.475 221.320 ;
        RECT 4.400 217.240 574.475 218.640 ;
        RECT 3.990 214.560 574.475 217.240 ;
        RECT 4.400 213.160 574.475 214.560 ;
        RECT 3.990 210.480 574.475 213.160 ;
        RECT 4.400 209.080 574.475 210.480 ;
        RECT 3.990 206.400 574.475 209.080 ;
        RECT 4.400 205.000 574.475 206.400 ;
        RECT 3.990 202.320 574.475 205.000 ;
        RECT 4.400 200.920 574.475 202.320 ;
        RECT 3.990 198.240 574.475 200.920 ;
        RECT 4.400 196.840 574.475 198.240 ;
        RECT 3.990 194.160 574.475 196.840 ;
        RECT 4.400 192.760 574.475 194.160 ;
        RECT 3.990 190.080 574.475 192.760 ;
        RECT 4.400 188.680 574.475 190.080 ;
        RECT 3.990 186.000 574.475 188.680 ;
        RECT 4.400 184.600 574.475 186.000 ;
        RECT 3.990 181.920 574.475 184.600 ;
        RECT 4.400 180.520 574.475 181.920 ;
        RECT 3.990 177.840 574.475 180.520 ;
        RECT 4.400 176.440 574.475 177.840 ;
        RECT 3.990 173.760 574.475 176.440 ;
        RECT 4.400 172.360 574.475 173.760 ;
        RECT 3.990 169.680 574.475 172.360 ;
        RECT 4.400 168.280 574.475 169.680 ;
        RECT 3.990 165.600 574.475 168.280 ;
        RECT 4.400 164.200 574.475 165.600 ;
        RECT 3.990 161.520 574.475 164.200 ;
        RECT 4.400 160.120 574.475 161.520 ;
        RECT 3.990 157.440 574.475 160.120 ;
        RECT 4.400 156.040 574.475 157.440 ;
        RECT 3.990 153.360 574.475 156.040 ;
        RECT 4.400 151.960 574.475 153.360 ;
        RECT 3.990 149.280 574.475 151.960 ;
        RECT 4.400 147.880 574.475 149.280 ;
        RECT 3.990 145.200 574.475 147.880 ;
        RECT 4.400 143.800 574.475 145.200 ;
        RECT 3.990 141.120 574.475 143.800 ;
        RECT 4.400 139.720 574.475 141.120 ;
        RECT 3.990 137.040 574.475 139.720 ;
        RECT 4.400 135.640 574.475 137.040 ;
        RECT 3.990 132.960 574.475 135.640 ;
        RECT 4.400 131.560 574.475 132.960 ;
        RECT 3.990 128.880 574.475 131.560 ;
        RECT 4.400 127.480 574.475 128.880 ;
        RECT 3.990 124.800 574.475 127.480 ;
        RECT 4.400 123.400 574.475 124.800 ;
        RECT 3.990 120.720 574.475 123.400 ;
        RECT 4.400 119.320 574.475 120.720 ;
        RECT 3.990 116.640 574.475 119.320 ;
        RECT 4.400 115.240 574.475 116.640 ;
        RECT 3.990 112.560 574.475 115.240 ;
        RECT 4.400 111.160 574.475 112.560 ;
        RECT 3.990 108.480 574.475 111.160 ;
        RECT 4.400 107.080 574.475 108.480 ;
        RECT 3.990 104.400 574.475 107.080 ;
        RECT 4.400 103.000 574.475 104.400 ;
        RECT 3.990 100.320 574.475 103.000 ;
        RECT 4.400 98.920 574.475 100.320 ;
        RECT 3.990 96.240 574.475 98.920 ;
        RECT 4.400 94.840 574.475 96.240 ;
        RECT 3.990 92.160 574.475 94.840 ;
        RECT 4.400 90.760 574.475 92.160 ;
        RECT 3.990 88.080 574.475 90.760 ;
        RECT 4.400 86.680 574.475 88.080 ;
        RECT 3.990 84.000 574.475 86.680 ;
        RECT 4.400 82.600 574.475 84.000 ;
        RECT 3.990 79.920 574.475 82.600 ;
        RECT 4.400 78.520 574.475 79.920 ;
        RECT 3.990 75.840 574.475 78.520 ;
        RECT 4.400 74.440 574.475 75.840 ;
        RECT 3.990 71.760 574.475 74.440 ;
        RECT 4.400 70.360 574.475 71.760 ;
        RECT 3.990 10.715 574.475 70.360 ;
      LAYER met4 ;
        RECT 19.615 59.335 20.640 559.465 ;
        RECT 23.040 59.335 97.440 559.465 ;
        RECT 99.840 59.335 174.240 559.465 ;
        RECT 176.640 59.335 251.040 559.465 ;
        RECT 253.440 59.335 327.840 559.465 ;
        RECT 330.240 59.335 404.640 559.465 ;
        RECT 407.040 59.335 481.440 559.465 ;
        RECT 483.840 59.335 558.145 559.465 ;
  END
END registerFile
END LIBRARY

